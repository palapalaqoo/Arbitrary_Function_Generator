`timescale	1ns/1ps

module	DECODE_DAC7821(DECODE_OUT, ADDR_IN, Clock)	;

output	[11:0]	DECODE_OUT	;
reg	[11:0]	DECODE_OUT	;

input	[25:0]	ADDR_IN	;
wire	[25:0]	ADDR_IN	;

input	Clock	;
wire	Clock	;


always	@(posedge	Clock)
	begin
		case(ADDR_IN)
		// A25A24.......................A3A2A1A0....................(A0 not used).....................
			26'b10_0000_0000_0000_0000_1010_0010 : DECODE_OUT <= 12'b0000_0000_0001	;		//DAC7821 MOD WAVE Value Enable................... 
			26'b10_0000_0000_0000_0000_1010_0100 : DECODE_OUT <= 12'b0000_0000_0010	;		//DAC7821 DC Offset Value Enable................... 
			26'b10_0000_0000_0000_0000_1010_0110 : DECODE_OUT <= 12'b0000_0000_0100	;		//DAC7821 Duty_S Value Enable................... 
			26'b10_0000_0000_0000_0000_1010_1000 : DECODE_OUT <= 12'b0000_0000_1000	;		//DAC7821 GAIN_V Value Enable................... 
			
			26'b10_0000_0000_0000_0000_1010_1010 : DECODE_OUT <= 12'b0000_0001_0000	;		//DAC7821 SQ_VL Value Enable...................
			26'b10_0000_0000_0000_0000_1010_1100 : DECODE_OUT <= 12'b0000_0010_0000	;		//DAC7821 SQ_VT Value Enable...................
			26'b10_0000_0000_0000_0000_1010_1110 : DECODE_OUT <= 12'b0000_0100_0000	;		//DAC7821 Spare Value Enable...................
			26'b10_0000_0000_0000_0000_1011_0000 : DECODE_OUT <= 12'b0000_1000_0000	;		//AM_Constants ..................
			
			26'b10_0000_0000_0000_0000_1011_0010 : DECODE_OUT <= 12'b0001_0000_0000	;		//Keypad Data Value Enable..................
			26'b10_0000_0000_0000_0000_1011_0100 : DECODE_OUT <= 12'b0010_0000_0000	;		//Reserved..................
			26'b10_0000_0000_0000_0000_1011_0110 : DECODE_OUT <= 12'b0100_0000_0000	;		//Reserved..................
			26'b10_0000_0000_0000_0000_1011_1000 : DECODE_OUT <= 12'b1000_0000_0000	;		//Reserved..................
			

			default : DECODE_OUT <= 12'b0000_0000_0000	;
		endcase
	end
	
endmodule


