//Look-Up Table for ROM of Version 4.....................
//The En pin must be connection to NRST..................


module	ROM_Table(Data_out, Addr_in, EN, Clock)	;

output	[15:0]	Data_out	;
reg	[15:0]	Data_out	;

input	[13:0]	Addr_in	;
wire	[13:0]	Addr_in	;

input	Clock	;
wire	Clock	;

input	EN	;
wire	EN	;


always	@(posedge	Clock)
	begin
		if ( EN == 1'b1 )
			case(Addr_in)
				/////////////////////////////////////////////////////////////////////////////////////////////
				//	posedge half-cycle of rise......
				14'b00000000000000: Data_out <= 16'h0000	;
				14'b00000000000001: Data_out <= 16'h000D	;
				14'b00000000000010: Data_out <= 16'h0019	;
				14'b00000000000011: Data_out <= 16'h0026	;
				14'b00000000000100: Data_out <= 16'h0032	;
				14'b00000000000101: Data_out <= 16'h003F	;
				14'b00000000000110: Data_out <= 16'h004B	;
				14'b00000000000111: Data_out <= 16'h0058	;
				14'b00000000001000: Data_out <= 16'h0065	;
				14'b00000000001001: Data_out <= 16'h0071	;
				14'b00000000001010: Data_out <= 16'h007E	;
				14'b00000000001011: Data_out <= 16'h008A	;
				14'b00000000001100: Data_out <= 16'h0097	;
				14'b00000000001101: Data_out <= 16'h00A3	;
				14'b00000000001110: Data_out <= 16'h00B0	;
				14'b00000000001111: Data_out <= 16'h00BD	;
				14'b00000000010000: Data_out <= 16'h00C9	;
				14'b00000000010001: Data_out <= 16'h00D6	;
				14'b00000000010010: Data_out <= 16'h00E2	;
				14'b00000000010011: Data_out <= 16'h00EF	;
				14'b00000000010100: Data_out <= 16'h00FB	;
				14'b00000000010101: Data_out <= 16'h0108	;
				14'b00000000010110: Data_out <= 16'h0115	;
				14'b00000000010111: Data_out <= 16'h0121	;
				14'b00000000011000: Data_out <= 16'h012E	;
				14'b00000000011001: Data_out <= 16'h013A	;
				14'b00000000011010: Data_out <= 16'h0147	;
				14'b00000000011011: Data_out <= 16'h0153	;
				14'b00000000011100: Data_out <= 16'h0160	;
				14'b00000000011101: Data_out <= 16'h016D	;
				14'b00000000011110: Data_out <= 16'h0179	;
				14'b00000000011111: Data_out <= 16'h0186	;
				14'b00000000100000: Data_out <= 16'h0192	;
				14'b00000000100001: Data_out <= 16'h019F	;
				14'b00000000100010: Data_out <= 16'h01AB	;
				14'b00000000100011: Data_out <= 16'h01B8	;
				14'b00000000100100: Data_out <= 16'h01C4	;
				14'b00000000100101: Data_out <= 16'h01D1	;
				14'b00000000100110: Data_out <= 16'h01DE	;
				14'b00000000100111: Data_out <= 16'h01EA	;
				14'b00000000101000: Data_out <= 16'h01F7	;
				14'b00000000101001: Data_out <= 16'h0203	;
				14'b00000000101010: Data_out <= 16'h0210	;
				14'b00000000101011: Data_out <= 16'h021C	;
				14'b00000000101100: Data_out <= 16'h0229	;
				14'b00000000101101: Data_out <= 16'h0236	;
				14'b00000000101110: Data_out <= 16'h0242	;
				14'b00000000101111: Data_out <= 16'h024F	;
				14'b00000000110000: Data_out <= 16'h025B	;
				14'b00000000110001: Data_out <= 16'h0268	;
				14'b00000000110010: Data_out <= 16'h0274	;
				14'b00000000110011: Data_out <= 16'h0281	;
				14'b00000000110100: Data_out <= 16'h028D	;
				14'b00000000110101: Data_out <= 16'h029A	;
				14'b00000000110110: Data_out <= 16'h02A7	;
				14'b00000000110111: Data_out <= 16'h02B3	;
				14'b00000000111000: Data_out <= 16'h02C0	;
				14'b00000000111001: Data_out <= 16'h02CC	;
				14'b00000000111010: Data_out <= 16'h02D9	;
				14'b00000000111011: Data_out <= 16'h02E5	;
				14'b00000000111100: Data_out <= 16'h02F2	;
				14'b00000000111101: Data_out <= 16'h02FF	;
				14'b00000000111110: Data_out <= 16'h030B	;
				14'b00000000111111: Data_out <= 16'h0318	;
				14'b00000001000000: Data_out <= 16'h0324	;
				14'b00000001000001: Data_out <= 16'h0331	;
				14'b00000001000010: Data_out <= 16'h033D	;
				14'b00000001000011: Data_out <= 16'h034A	;
				14'b00000001000100: Data_out <= 16'h0356	;
				14'b00000001000101: Data_out <= 16'h0363	;
				14'b00000001000110: Data_out <= 16'h0370	;
				14'b00000001000111: Data_out <= 16'h037C	;
				14'b00000001001000: Data_out <= 16'h0389	;
				14'b00000001001001: Data_out <= 16'h0395	;
				14'b00000001001010: Data_out <= 16'h03A2	;
				14'b00000001001011: Data_out <= 16'h03AE	;
				14'b00000001001100: Data_out <= 16'h03BB	;
				14'b00000001001101: Data_out <= 16'h03C8	;
				14'b00000001001110: Data_out <= 16'h03D4	;
				14'b00000001001111: Data_out <= 16'h03E1	;
				14'b00000001010000: Data_out <= 16'h03ED	;
				14'b00000001010001: Data_out <= 16'h03FA	;
				14'b00000001010010: Data_out <= 16'h0406	;
				14'b00000001010011: Data_out <= 16'h0413	;
				14'b00000001010100: Data_out <= 16'h041F	;
				14'b00000001010101: Data_out <= 16'h042C	;
				14'b00000001010110: Data_out <= 16'h0439	;
				14'b00000001010111: Data_out <= 16'h0445	;
				14'b00000001011000: Data_out <= 16'h0452	;
				14'b00000001011001: Data_out <= 16'h045E	;
				14'b00000001011010: Data_out <= 16'h046B	;
				14'b00000001011011: Data_out <= 16'h0477	;
				14'b00000001011100: Data_out <= 16'h0484	;
				14'b00000001011101: Data_out <= 16'h0490	;
				14'b00000001011110: Data_out <= 16'h049D	;
				14'b00000001011111: Data_out <= 16'h04AA	;
				14'b00000001100000: Data_out <= 16'h04B6	;
				14'b00000001100001: Data_out <= 16'h04C3	;
				14'b00000001100010: Data_out <= 16'h04CF	;
				14'b00000001100011: Data_out <= 16'h04DC	;
				14'b00000001100100: Data_out <= 16'h04E8	;
				14'b00000001100101: Data_out <= 16'h04F5	;
				14'b00000001100110: Data_out <= 16'h0502	;
				14'b00000001100111: Data_out <= 16'h050E	;
				14'b00000001101000: Data_out <= 16'h051B	;
				14'b00000001101001: Data_out <= 16'h0527	;
				14'b00000001101010: Data_out <= 16'h0534	;
				14'b00000001101011: Data_out <= 16'h0540	;
				14'b00000001101100: Data_out <= 16'h054D	;
				14'b00000001101101: Data_out <= 16'h0559	;
				14'b00000001101110: Data_out <= 16'h0566	;
				14'b00000001101111: Data_out <= 16'h0573	;
				14'b00000001110000: Data_out <= 16'h057F	;
				14'b00000001110001: Data_out <= 16'h058C	;
				14'b00000001110010: Data_out <= 16'h0598	;
				14'b00000001110011: Data_out <= 16'h05A5	;
				14'b00000001110100: Data_out <= 16'h05B1	;
				14'b00000001110101: Data_out <= 16'h05BE	;
				14'b00000001110110: Data_out <= 16'h05CA	;
				14'b00000001110111: Data_out <= 16'h05D7	;
				14'b00000001111000: Data_out <= 16'h05E3	;
				14'b00000001111001: Data_out <= 16'h05F0	;
				14'b00000001111010: Data_out <= 16'h05FD	;
				14'b00000001111011: Data_out <= 16'h0609	;
				14'b00000001111100: Data_out <= 16'h0616	;
				14'b00000001111101: Data_out <= 16'h0622	;
				14'b00000001111110: Data_out <= 16'h062F	;
				14'b00000001111111: Data_out <= 16'h063B	;
				14'b00000010000000: Data_out <= 16'h0648	;
				14'b00000010000001: Data_out <= 16'h0654	;
				14'b00000010000010: Data_out <= 16'h0661	;
				14'b00000010000011: Data_out <= 16'h066E	;
				14'b00000010000100: Data_out <= 16'h067A	;
				14'b00000010000101: Data_out <= 16'h0687	;
				14'b00000010000110: Data_out <= 16'h0693	;
				14'b00000010000111: Data_out <= 16'h06A0	;
				14'b00000010001000: Data_out <= 16'h06AC	;
				14'b00000010001001: Data_out <= 16'h06B9	;
				14'b00000010001010: Data_out <= 16'h06C5	;
				14'b00000010001011: Data_out <= 16'h06D2	;
				14'b00000010001100: Data_out <= 16'h06DE	;
				14'b00000010001101: Data_out <= 16'h06EB	;
				14'b00000010001110: Data_out <= 16'h06F8	;
				14'b00000010001111: Data_out <= 16'h0704	;
				14'b00000010010000: Data_out <= 16'h0711	;
				14'b00000010010001: Data_out <= 16'h071D	;
				14'b00000010010010: Data_out <= 16'h072A	;
				14'b00000010010011: Data_out <= 16'h0736	;
				14'b00000010010100: Data_out <= 16'h0743	;
				14'b00000010010101: Data_out <= 16'h074F	;
				14'b00000010010110: Data_out <= 16'h075C	;
				14'b00000010010111: Data_out <= 16'h0769	;
				14'b00000010011000: Data_out <= 16'h0775	;
				14'b00000010011001: Data_out <= 16'h0782	;
				14'b00000010011010: Data_out <= 16'h078E	;
				14'b00000010011011: Data_out <= 16'h079B	;
				14'b00000010011100: Data_out <= 16'h07A7	;
				14'b00000010011101: Data_out <= 16'h07B4	;
				14'b00000010011110: Data_out <= 16'h07C0	;
				14'b00000010011111: Data_out <= 16'h07CD	;
				14'b00000010100000: Data_out <= 16'h07D9	;
				14'b00000010100001: Data_out <= 16'h07E6	;
				14'b00000010100010: Data_out <= 16'h07F2	;
				14'b00000010100011: Data_out <= 16'h07FF	;
				14'b00000010100100: Data_out <= 16'h080C	;
				14'b00000010100101: Data_out <= 16'h0818	;
				14'b00000010100110: Data_out <= 16'h0825	;
				14'b00000010100111: Data_out <= 16'h0831	;
				14'b00000010101000: Data_out <= 16'h083E	;
				14'b00000010101001: Data_out <= 16'h084A	;
				14'b00000010101010: Data_out <= 16'h0857	;
				14'b00000010101011: Data_out <= 16'h0863	;
				14'b00000010101100: Data_out <= 16'h0870	;
				14'b00000010101101: Data_out <= 16'h087C	;
				14'b00000010101110: Data_out <= 16'h0889	;
				14'b00000010101111: Data_out <= 16'h0895	;
				14'b00000010110000: Data_out <= 16'h08A2	;
				14'b00000010110001: Data_out <= 16'h08AF	;
				14'b00000010110010: Data_out <= 16'h08BB	;
				14'b00000010110011: Data_out <= 16'h08C8	;
				14'b00000010110100: Data_out <= 16'h08D4	;
				14'b00000010110101: Data_out <= 16'h08E1	;
				14'b00000010110110: Data_out <= 16'h08ED	;
				14'b00000010110111: Data_out <= 16'h08FA	;
				14'b00000010111000: Data_out <= 16'h0906	;
				14'b00000010111001: Data_out <= 16'h0913	;
				14'b00000010111010: Data_out <= 16'h091F	;
				14'b00000010111011: Data_out <= 16'h092C	;
				14'b00000010111100: Data_out <= 16'h0938	;
				14'b00000010111101: Data_out <= 16'h0945	;
				14'b00000010111110: Data_out <= 16'h0952	;
				14'b00000010111111: Data_out <= 16'h095E	;
				14'b00000011000000: Data_out <= 16'h096B	;
				14'b00000011000001: Data_out <= 16'h0977	;
				14'b00000011000010: Data_out <= 16'h0984	;
				14'b00000011000011: Data_out <= 16'h0990	;
				14'b00000011000100: Data_out <= 16'h099D	;
				14'b00000011000101: Data_out <= 16'h09A9	;
				14'b00000011000110: Data_out <= 16'h09B6	;
				14'b00000011000111: Data_out <= 16'h09C2	;
				14'b00000011001000: Data_out <= 16'h09CF	;
				14'b00000011001001: Data_out <= 16'h09DB	;
				14'b00000011001010: Data_out <= 16'h09E8	;
				14'b00000011001011: Data_out <= 16'h09F4	;
				14'b00000011001100: Data_out <= 16'h0A01	;
				14'b00000011001101: Data_out <= 16'h0A0D	;
				14'b00000011001110: Data_out <= 16'h0A1A	;
				14'b00000011001111: Data_out <= 16'h0A27	;
				14'b00000011010000: Data_out <= 16'h0A33	;
				14'b00000011010001: Data_out <= 16'h0A40	;
				14'b00000011010010: Data_out <= 16'h0A4C	;
				14'b00000011010011: Data_out <= 16'h0A59	;
				14'b00000011010100: Data_out <= 16'h0A65	;
				14'b00000011010101: Data_out <= 16'h0A72	;
				14'b00000011010110: Data_out <= 16'h0A7E	;
				14'b00000011010111: Data_out <= 16'h0A8B	;
				14'b00000011011000: Data_out <= 16'h0A97	;
				14'b00000011011001: Data_out <= 16'h0AA4	;
				14'b00000011011010: Data_out <= 16'h0AB0	;
				14'b00000011011011: Data_out <= 16'h0ABD	;
				14'b00000011011100: Data_out <= 16'h0AC9	;
				14'b00000011011101: Data_out <= 16'h0AD6	;
				14'b00000011011110: Data_out <= 16'h0AE2	;
				14'b00000011011111: Data_out <= 16'h0AEF	;
				14'b00000011100000: Data_out <= 16'h0AFB	;
				14'b00000011100001: Data_out <= 16'h0B08	;
				14'b00000011100010: Data_out <= 16'h0B14	;
				14'b00000011100011: Data_out <= 16'h0B21	;
				14'b00000011100100: Data_out <= 16'h0B2D	;
				14'b00000011100101: Data_out <= 16'h0B3A	;
				14'b00000011100110: Data_out <= 16'h0B47	;
				14'b00000011100111: Data_out <= 16'h0B53	;
				14'b00000011101000: Data_out <= 16'h0B60	;
				14'b00000011101001: Data_out <= 16'h0B6C	;
				14'b00000011101010: Data_out <= 16'h0B79	;
				14'b00000011101011: Data_out <= 16'h0B85	;
				14'b00000011101100: Data_out <= 16'h0B92	;
				14'b00000011101101: Data_out <= 16'h0B9E	;
				14'b00000011101110: Data_out <= 16'h0BAB	;
				14'b00000011101111: Data_out <= 16'h0BB7	;
				14'b00000011110000: Data_out <= 16'h0BC4	;
				14'b00000011110001: Data_out <= 16'h0BD0	;
				14'b00000011110010: Data_out <= 16'h0BDD	;
				14'b00000011110011: Data_out <= 16'h0BE9	;
				14'b00000011110100: Data_out <= 16'h0BF6	;
				14'b00000011110101: Data_out <= 16'h0C02	;
				14'b00000011110110: Data_out <= 16'h0C0F	;
				14'b00000011110111: Data_out <= 16'h0C1B	;
				14'b00000011111000: Data_out <= 16'h0C28	;
				14'b00000011111001: Data_out <= 16'h0C34	;
				14'b00000011111010: Data_out <= 16'h0C41	;
				14'b00000011111011: Data_out <= 16'h0C4D	;
				14'b00000011111100: Data_out <= 16'h0C5A	;
				14'b00000011111101: Data_out <= 16'h0C66	;
				14'b00000011111110: Data_out <= 16'h0C73	;
				14'b00000011111111: Data_out <= 16'h0C7F	;
				14'b00000100000000: Data_out <= 16'h0C8C	;
				14'b00000100000001: Data_out <= 16'h0C98	;
				14'b00000100000010: Data_out <= 16'h0CA5	;
				14'b00000100000011: Data_out <= 16'h0CB1	;
				14'b00000100000100: Data_out <= 16'h0CBE	;
				14'b00000100000101: Data_out <= 16'h0CCA	;
				14'b00000100000110: Data_out <= 16'h0CD7	;
				14'b00000100000111: Data_out <= 16'h0CE3	;
				14'b00000100001000: Data_out <= 16'h0CF0	;
				14'b00000100001001: Data_out <= 16'h0CFC	;
				14'b00000100001010: Data_out <= 16'h0D09	;
				14'b00000100001011: Data_out <= 16'h0D15	;
				14'b00000100001100: Data_out <= 16'h0D22	;
				14'b00000100001101: Data_out <= 16'h0D2E	;
				14'b00000100001110: Data_out <= 16'h0D3B	;
				14'b00000100001111: Data_out <= 16'h0D47	;
				14'b00000100010000: Data_out <= 16'h0D54	;
				14'b00000100010001: Data_out <= 16'h0D60	;
				14'b00000100010010: Data_out <= 16'h0D6D	;
				14'b00000100010011: Data_out <= 16'h0D79	;
				14'b00000100010100: Data_out <= 16'h0D86	;
				14'b00000100010101: Data_out <= 16'h0D92	;
				14'b00000100010110: Data_out <= 16'h0D9F	;
				14'b00000100010111: Data_out <= 16'h0DAB	;
				14'b00000100011000: Data_out <= 16'h0DB8	;
				14'b00000100011001: Data_out <= 16'h0DC4	;
				14'b00000100011010: Data_out <= 16'h0DD1	;
				14'b00000100011011: Data_out <= 16'h0DDD	;
				14'b00000100011100: Data_out <= 16'h0DEA	;
				14'b00000100011101: Data_out <= 16'h0DF6	;
				14'b00000100011110: Data_out <= 16'h0E03	;
				14'b00000100011111: Data_out <= 16'h0E0F	;
				14'b00000100100000: Data_out <= 16'h0E1C	;
				14'b00000100100001: Data_out <= 16'h0E28	;
				14'b00000100100010: Data_out <= 16'h0E35	;
				14'b00000100100011: Data_out <= 16'h0E41	;
				14'b00000100100100: Data_out <= 16'h0E4E	;
				14'b00000100100101: Data_out <= 16'h0E5A	;
				14'b00000100100110: Data_out <= 16'h0E67	;
				14'b00000100100111: Data_out <= 16'h0E73	;
				14'b00000100101000: Data_out <= 16'h0E80	;
				14'b00000100101001: Data_out <= 16'h0E8C	;
				14'b00000100101010: Data_out <= 16'h0E99	;
				14'b00000100101011: Data_out <= 16'h0EA5	;
				14'b00000100101100: Data_out <= 16'h0EB2	;
				14'b00000100101101: Data_out <= 16'h0EBE	;
				14'b00000100101110: Data_out <= 16'h0ECB	;
				14'b00000100101111: Data_out <= 16'h0ED7	;
				14'b00000100110000: Data_out <= 16'h0EE4	;
				14'b00000100110001: Data_out <= 16'h0EF0	;
				14'b00000100110010: Data_out <= 16'h0EFC	;
				14'b00000100110011: Data_out <= 16'h0F09	;
				14'b00000100110100: Data_out <= 16'h0F15	;
				14'b00000100110101: Data_out <= 16'h0F22	;
				14'b00000100110110: Data_out <= 16'h0F2E	;
				14'b00000100110111: Data_out <= 16'h0F3B	;
				14'b00000100111000: Data_out <= 16'h0F47	;
				14'b00000100111001: Data_out <= 16'h0F54	;
				14'b00000100111010: Data_out <= 16'h0F60	;
				14'b00000100111011: Data_out <= 16'h0F6D	;
				14'b00000100111100: Data_out <= 16'h0F79	;
				14'b00000100111101: Data_out <= 16'h0F86	;
				14'b00000100111110: Data_out <= 16'h0F92	;
				14'b00000100111111: Data_out <= 16'h0F9F	;
				14'b00000101000000: Data_out <= 16'h0FAB	;
				14'b00000101000001: Data_out <= 16'h0FB8	;
				14'b00000101000010: Data_out <= 16'h0FC4	;
				14'b00000101000011: Data_out <= 16'h0FD1	;
				14'b00000101000100: Data_out <= 16'h0FDD	;
				14'b00000101000101: Data_out <= 16'h0FE9	;
				14'b00000101000110: Data_out <= 16'h0FF6	;
				14'b00000101000111: Data_out <= 16'h1002	;
				14'b00000101001000: Data_out <= 16'h100F	;
				14'b00000101001001: Data_out <= 16'h101B	;
				14'b00000101001010: Data_out <= 16'h1028	;
				14'b00000101001011: Data_out <= 16'h1034	;
				14'b00000101001100: Data_out <= 16'h1041	;
				14'b00000101001101: Data_out <= 16'h104D	;
				14'b00000101001110: Data_out <= 16'h105A	;
				14'b00000101001111: Data_out <= 16'h1066	;
				14'b00000101010000: Data_out <= 16'h1073	;
				14'b00000101010001: Data_out <= 16'h107F	;
				14'b00000101010010: Data_out <= 16'h108C	;
				14'b00000101010011: Data_out <= 16'h1098	;
				14'b00000101010100: Data_out <= 16'h10A4	;
				14'b00000101010101: Data_out <= 16'h10B1	;
				14'b00000101010110: Data_out <= 16'h10BD	;
				14'b00000101010111: Data_out <= 16'h10CA	;
				14'b00000101011000: Data_out <= 16'h10D6	;
				14'b00000101011001: Data_out <= 16'h10E3	;
				14'b00000101011010: Data_out <= 16'h10EF	;
				14'b00000101011011: Data_out <= 16'h10FC	;
				14'b00000101011100: Data_out <= 16'h1108	;
				14'b00000101011101: Data_out <= 16'h1115	;
				14'b00000101011110: Data_out <= 16'h1121	;
				14'b00000101011111: Data_out <= 16'h112D	;
				14'b00000101100000: Data_out <= 16'h113A	;
				14'b00000101100001: Data_out <= 16'h1146	;
				14'b00000101100010: Data_out <= 16'h1153	;
				14'b00000101100011: Data_out <= 16'h115F	;
				14'b00000101100100: Data_out <= 16'h116C	;
				14'b00000101100101: Data_out <= 16'h1178	;
				14'b00000101100110: Data_out <= 16'h1185	;
				14'b00000101100111: Data_out <= 16'h1191	;
				14'b00000101101000: Data_out <= 16'h119D	;
				14'b00000101101001: Data_out <= 16'h11AA	;
				14'b00000101101010: Data_out <= 16'h11B6	;
				14'b00000101101011: Data_out <= 16'h11C3	;
				14'b00000101101100: Data_out <= 16'h11CF	;
				14'b00000101101101: Data_out <= 16'h11DC	;
				14'b00000101101110: Data_out <= 16'h11E8	;
				14'b00000101101111: Data_out <= 16'h11F5	;
				14'b00000101110000: Data_out <= 16'h1201	;
				14'b00000101110001: Data_out <= 16'h120D	;
				14'b00000101110010: Data_out <= 16'h121A	;
				14'b00000101110011: Data_out <= 16'h1226	;
				14'b00000101110100: Data_out <= 16'h1233	;
				14'b00000101110101: Data_out <= 16'h123F	;
				14'b00000101110110: Data_out <= 16'h124C	;
				14'b00000101110111: Data_out <= 16'h1258	;
				14'b00000101111000: Data_out <= 16'h1265	;
				14'b00000101111001: Data_out <= 16'h1271	;
				14'b00000101111010: Data_out <= 16'h127D	;
				14'b00000101111011: Data_out <= 16'h128A	;
				14'b00000101111100: Data_out <= 16'h1296	;
				14'b00000101111101: Data_out <= 16'h12A3	;
				14'b00000101111110: Data_out <= 16'h12AF	;
				14'b00000101111111: Data_out <= 16'h12BC	;
				14'b00000110000000: Data_out <= 16'h12C8	;
				14'b00000110000001: Data_out <= 16'h12D4	;
				14'b00000110000010: Data_out <= 16'h12E1	;
				14'b00000110000011: Data_out <= 16'h12ED	;
				14'b00000110000100: Data_out <= 16'h12FA	;
				14'b00000110000101: Data_out <= 16'h1306	;
				14'b00000110000110: Data_out <= 16'h1313	;
				14'b00000110000111: Data_out <= 16'h131F	;
				14'b00000110001000: Data_out <= 16'h132B	;
				14'b00000110001001: Data_out <= 16'h1338	;
				14'b00000110001010: Data_out <= 16'h1344	;
				14'b00000110001011: Data_out <= 16'h1351	;
				14'b00000110001100: Data_out <= 16'h135D	;
				14'b00000110001101: Data_out <= 16'h136A	;
				14'b00000110001110: Data_out <= 16'h1376	;
				14'b00000110001111: Data_out <= 16'h1382	;
				14'b00000110010000: Data_out <= 16'h138F	;
				14'b00000110010001: Data_out <= 16'h139B	;
				14'b00000110010010: Data_out <= 16'h13A8	;
				14'b00000110010011: Data_out <= 16'h13B4	;
				14'b00000110010100: Data_out <= 16'h13C0	;
				14'b00000110010101: Data_out <= 16'h13CD	;
				14'b00000110010110: Data_out <= 16'h13D9	;
				14'b00000110010111: Data_out <= 16'h13E6	;
				14'b00000110011000: Data_out <= 16'h13F2	;
				14'b00000110011001: Data_out <= 16'h13FF	;
				14'b00000110011010: Data_out <= 16'h140B	;
				14'b00000110011011: Data_out <= 16'h1417	;
				14'b00000110011100: Data_out <= 16'h1424	;
				14'b00000110011101: Data_out <= 16'h1430	;
				14'b00000110011110: Data_out <= 16'h143D	;
				14'b00000110011111: Data_out <= 16'h1449	;
				14'b00000110100000: Data_out <= 16'h1455	;
				14'b00000110100001: Data_out <= 16'h1462	;
				14'b00000110100010: Data_out <= 16'h146E	;
				14'b00000110100011: Data_out <= 16'h147B	;
				14'b00000110100100: Data_out <= 16'h1487	;
				14'b00000110100101: Data_out <= 16'h1493	;
				14'b00000110100110: Data_out <= 16'h14A0	;
				14'b00000110100111: Data_out <= 16'h14AC	;
				14'b00000110101000: Data_out <= 16'h14B9	;
				14'b00000110101001: Data_out <= 16'h14C5	;
				14'b00000110101010: Data_out <= 16'h14D1	;
				14'b00000110101011: Data_out <= 16'h14DE	;
				14'b00000110101100: Data_out <= 16'h14EA	;
				14'b00000110101101: Data_out <= 16'h14F7	;
				14'b00000110101110: Data_out <= 16'h1503	;
				14'b00000110101111: Data_out <= 16'h150F	;
				14'b00000110110000: Data_out <= 16'h151C	;
				14'b00000110110001: Data_out <= 16'h1528	;
				14'b00000110110010: Data_out <= 16'h1535	;
				14'b00000110110011: Data_out <= 16'h1541	;
				14'b00000110110100: Data_out <= 16'h154D	;
				14'b00000110110101: Data_out <= 16'h155A	;
				14'b00000110110110: Data_out <= 16'h1566	;
				14'b00000110110111: Data_out <= 16'h1573	;
				14'b00000110111000: Data_out <= 16'h157F	;
				14'b00000110111001: Data_out <= 16'h158B	;
				14'b00000110111010: Data_out <= 16'h1598	;
				14'b00000110111011: Data_out <= 16'h15A4	;
				14'b00000110111100: Data_out <= 16'h15B0	;
				14'b00000110111101: Data_out <= 16'h15BD	;
				14'b00000110111110: Data_out <= 16'h15C9	;
				14'b00000110111111: Data_out <= 16'h15D6	;
				14'b00000111000000: Data_out <= 16'h15E2	;
				14'b00000111000001: Data_out <= 16'h15EE	;
				14'b00000111000010: Data_out <= 16'h15FB	;
				14'b00000111000011: Data_out <= 16'h1607	;
				14'b00000111000100: Data_out <= 16'h1614	;
				14'b00000111000101: Data_out <= 16'h1620	;
				14'b00000111000110: Data_out <= 16'h162C	;
				14'b00000111000111: Data_out <= 16'h1639	;
				14'b00000111001000: Data_out <= 16'h1645	;
				14'b00000111001001: Data_out <= 16'h1651	;
				14'b00000111001010: Data_out <= 16'h165E	;
				14'b00000111001011: Data_out <= 16'h166A	;
				14'b00000111001100: Data_out <= 16'h1677	;
				14'b00000111001101: Data_out <= 16'h1683	;
				14'b00000111001110: Data_out <= 16'h168F	;
				14'b00000111001111: Data_out <= 16'h169C	;
				14'b00000111010000: Data_out <= 16'h16A8	;
				14'b00000111010001: Data_out <= 16'h16B4	;
				14'b00000111010010: Data_out <= 16'h16C1	;
				14'b00000111010011: Data_out <= 16'h16CD	;
				14'b00000111010100: Data_out <= 16'h16D9	;
				14'b00000111010101: Data_out <= 16'h16E6	;
				14'b00000111010110: Data_out <= 16'h16F2	;
				14'b00000111010111: Data_out <= 16'h16FF	;
				14'b00000111011000: Data_out <= 16'h170B	;
				14'b00000111011001: Data_out <= 16'h1717	;
				14'b00000111011010: Data_out <= 16'h1724	;
				14'b00000111011011: Data_out <= 16'h1730	;
				14'b00000111011100: Data_out <= 16'h173C	;
				14'b00000111011101: Data_out <= 16'h1749	;
				14'b00000111011110: Data_out <= 16'h1755	;
				14'b00000111011111: Data_out <= 16'h1761	;
				14'b00000111100000: Data_out <= 16'h176E	;
				14'b00000111100001: Data_out <= 16'h177A	;
				14'b00000111100010: Data_out <= 16'h1786	;
				14'b00000111100011: Data_out <= 16'h1793	;
				14'b00000111100100: Data_out <= 16'h179F	;
				14'b00000111100101: Data_out <= 16'h17AC	;
				14'b00000111100110: Data_out <= 16'h17B8	;
				14'b00000111100111: Data_out <= 16'h17C4	;
				14'b00000111101000: Data_out <= 16'h17D1	;
				14'b00000111101001: Data_out <= 16'h17DD	;
				14'b00000111101010: Data_out <= 16'h17E9	;
				14'b00000111101011: Data_out <= 16'h17F6	;
				14'b00000111101100: Data_out <= 16'h1802	;
				14'b00000111101101: Data_out <= 16'h180E	;
				14'b00000111101110: Data_out <= 16'h181B	;
				14'b00000111101111: Data_out <= 16'h1827	;
				14'b00000111110000: Data_out <= 16'h1833	;
				14'b00000111110001: Data_out <= 16'h1840	;
				14'b00000111110010: Data_out <= 16'h184C	;
				14'b00000111110011: Data_out <= 16'h1858	;
				14'b00000111110100: Data_out <= 16'h1865	;
				14'b00000111110101: Data_out <= 16'h1871	;
				14'b00000111110110: Data_out <= 16'h187D	;
				14'b00000111110111: Data_out <= 16'h188A	;
				14'b00000111111000: Data_out <= 16'h1896	;
				14'b00000111111001: Data_out <= 16'h18A2	;
				14'b00000111111010: Data_out <= 16'h18AF	;
				14'b00000111111011: Data_out <= 16'h18BB	;
				14'b00000111111100: Data_out <= 16'h18C7	;
				14'b00000111111101: Data_out <= 16'h18D4	;
				14'b00000111111110: Data_out <= 16'h18E0	;
				14'b00000111111111: Data_out <= 16'h18EC	;
				14'b00001000000000: Data_out <= 16'h18F9	;
				14'b00001000000001: Data_out <= 16'h1905	;
				14'b00001000000010: Data_out <= 16'h1911	;
				14'b00001000000011: Data_out <= 16'h191E	;
				14'b00001000000100: Data_out <= 16'h192A	;
				14'b00001000000101: Data_out <= 16'h1936	;
				14'b00001000000110: Data_out <= 16'h1943	;
				14'b00001000000111: Data_out <= 16'h194F	;
				14'b00001000001000: Data_out <= 16'h195B	;
				14'b00001000001001: Data_out <= 16'h1968	;
				14'b00001000001010: Data_out <= 16'h1974	;
				14'b00001000001011: Data_out <= 16'h1980	;
				14'b00001000001100: Data_out <= 16'h198C	;
				14'b00001000001101: Data_out <= 16'h1999	;
				14'b00001000001110: Data_out <= 16'h19A5	;
				14'b00001000001111: Data_out <= 16'h19B1	;
				14'b00001000010000: Data_out <= 16'h19BE	;
				14'b00001000010001: Data_out <= 16'h19CA	;
				14'b00001000010010: Data_out <= 16'h19D6	;
				14'b00001000010011: Data_out <= 16'h19E3	;
				14'b00001000010100: Data_out <= 16'h19EF	;
				14'b00001000010101: Data_out <= 16'h19FB	;
				14'b00001000010110: Data_out <= 16'h1A08	;
				14'b00001000010111: Data_out <= 16'h1A14	;
				14'b00001000011000: Data_out <= 16'h1A20	;
				14'b00001000011001: Data_out <= 16'h1A2C	;
				14'b00001000011010: Data_out <= 16'h1A39	;
				14'b00001000011011: Data_out <= 16'h1A45	;
				14'b00001000011100: Data_out <= 16'h1A51	;
				14'b00001000011101: Data_out <= 16'h1A5E	;
				14'b00001000011110: Data_out <= 16'h1A6A	;
				14'b00001000011111: Data_out <= 16'h1A76	;
				14'b00001000100000: Data_out <= 16'h1A83	;
				14'b00001000100001: Data_out <= 16'h1A8F	;
				14'b00001000100010: Data_out <= 16'h1A9B	;
				14'b00001000100011: Data_out <= 16'h1AA7	;
				14'b00001000100100: Data_out <= 16'h1AB4	;
				14'b00001000100101: Data_out <= 16'h1AC0	;
				14'b00001000100110: Data_out <= 16'h1ACC	;
				14'b00001000100111: Data_out <= 16'h1AD9	;
				14'b00001000101000: Data_out <= 16'h1AE5	;
				14'b00001000101001: Data_out <= 16'h1AF1	;
				14'b00001000101010: Data_out <= 16'h1AFD	;
				14'b00001000101011: Data_out <= 16'h1B0A	;
				14'b00001000101100: Data_out <= 16'h1B16	;
				14'b00001000101101: Data_out <= 16'h1B22	;
				14'b00001000101110: Data_out <= 16'h1B2F	;
				14'b00001000101111: Data_out <= 16'h1B3B	;
				14'b00001000110000: Data_out <= 16'h1B47	;
				14'b00001000110001: Data_out <= 16'h1B53	;
				14'b00001000110010: Data_out <= 16'h1B60	;
				14'b00001000110011: Data_out <= 16'h1B6C	;
				14'b00001000110100: Data_out <= 16'h1B78	;
				14'b00001000110101: Data_out <= 16'h1B84	;
				14'b00001000110110: Data_out <= 16'h1B91	;
				14'b00001000110111: Data_out <= 16'h1B9D	;
				14'b00001000111000: Data_out <= 16'h1BA9	;
				14'b00001000111001: Data_out <= 16'h1BB6	;
				14'b00001000111010: Data_out <= 16'h1BC2	;
				14'b00001000111011: Data_out <= 16'h1BCE	;
				14'b00001000111100: Data_out <= 16'h1BDA	;
				14'b00001000111101: Data_out <= 16'h1BE7	;
				14'b00001000111110: Data_out <= 16'h1BF3	;
				14'b00001000111111: Data_out <= 16'h1BFF	;
				14'b00001001000000: Data_out <= 16'h1C0B	;
				14'b00001001000001: Data_out <= 16'h1C18	;
				14'b00001001000010: Data_out <= 16'h1C24	;
				14'b00001001000011: Data_out <= 16'h1C30	;
				14'b00001001000100: Data_out <= 16'h1C3C	;
				14'b00001001000101: Data_out <= 16'h1C49	;
				14'b00001001000110: Data_out <= 16'h1C55	;
				14'b00001001000111: Data_out <= 16'h1C61	;
				14'b00001001001000: Data_out <= 16'h1C6D	;
				14'b00001001001001: Data_out <= 16'h1C7A	;
				14'b00001001001010: Data_out <= 16'h1C86	;
				14'b00001001001011: Data_out <= 16'h1C92	;
				14'b00001001001100: Data_out <= 16'h1C9E	;
				14'b00001001001101: Data_out <= 16'h1CAB	;
				14'b00001001001110: Data_out <= 16'h1CB7	;
				14'b00001001001111: Data_out <= 16'h1CC3	;
				14'b00001001010000: Data_out <= 16'h1CCF	;
				14'b00001001010001: Data_out <= 16'h1CDC	;
				14'b00001001010010: Data_out <= 16'h1CE8	;
				14'b00001001010011: Data_out <= 16'h1CF4	;
				14'b00001001010100: Data_out <= 16'h1D00	;
				14'b00001001010101: Data_out <= 16'h1D0D	;
				14'b00001001010110: Data_out <= 16'h1D19	;
				14'b00001001010111: Data_out <= 16'h1D25	;
				14'b00001001011000: Data_out <= 16'h1D31	;
				14'b00001001011001: Data_out <= 16'h1D3E	;
				14'b00001001011010: Data_out <= 16'h1D4A	;
				14'b00001001011011: Data_out <= 16'h1D56	;
				14'b00001001011100: Data_out <= 16'h1D62	;
				14'b00001001011101: Data_out <= 16'h1D6E	;
				14'b00001001011110: Data_out <= 16'h1D7B	;
				14'b00001001011111: Data_out <= 16'h1D87	;
				14'b00001001100000: Data_out <= 16'h1D93	;
				14'b00001001100001: Data_out <= 16'h1D9F	;
				14'b00001001100010: Data_out <= 16'h1DAC	;
				14'b00001001100011: Data_out <= 16'h1DB8	;
				14'b00001001100100: Data_out <= 16'h1DC4	;
				14'b00001001100101: Data_out <= 16'h1DD0	;
				14'b00001001100110: Data_out <= 16'h1DDD	;
				14'b00001001100111: Data_out <= 16'h1DE9	;
				14'b00001001101000: Data_out <= 16'h1DF5	;
				14'b00001001101001: Data_out <= 16'h1E01	;
				14'b00001001101010: Data_out <= 16'h1E0D	;
				14'b00001001101011: Data_out <= 16'h1E1A	;
				14'b00001001101100: Data_out <= 16'h1E26	;
				14'b00001001101101: Data_out <= 16'h1E32	;
				14'b00001001101110: Data_out <= 16'h1E3E	;
				14'b00001001101111: Data_out <= 16'h1E4A	;
				14'b00001001110000: Data_out <= 16'h1E57	;
				14'b00001001110001: Data_out <= 16'h1E63	;
				14'b00001001110010: Data_out <= 16'h1E6F	;
				14'b00001001110011: Data_out <= 16'h1E7B	;
				14'b00001001110100: Data_out <= 16'h1E87	;
				14'b00001001110101: Data_out <= 16'h1E94	;
				14'b00001001110110: Data_out <= 16'h1EA0	;
				14'b00001001110111: Data_out <= 16'h1EAC	;
				14'b00001001111000: Data_out <= 16'h1EB8	;
				14'b00001001111001: Data_out <= 16'h1EC4	;
				14'b00001001111010: Data_out <= 16'h1ED1	;
				14'b00001001111011: Data_out <= 16'h1EDD	;
				14'b00001001111100: Data_out <= 16'h1EE9	;
				14'b00001001111101: Data_out <= 16'h1EF5	;
				14'b00001001111110: Data_out <= 16'h1F01	;
				14'b00001001111111: Data_out <= 16'h1F0E	;
				14'b00001010000000: Data_out <= 16'h1F1A	;
				14'b00001010000001: Data_out <= 16'h1F26	;
				14'b00001010000010: Data_out <= 16'h1F32	;
				14'b00001010000011: Data_out <= 16'h1F3E	;
				14'b00001010000100: Data_out <= 16'h1F4B	;
				14'b00001010000101: Data_out <= 16'h1F57	;
				14'b00001010000110: Data_out <= 16'h1F63	;
				14'b00001010000111: Data_out <= 16'h1F6F	;
				14'b00001010001000: Data_out <= 16'h1F7B	;
				14'b00001010001001: Data_out <= 16'h1F87	;
				14'b00001010001010: Data_out <= 16'h1F94	;
				14'b00001010001011: Data_out <= 16'h1FA0	;
				14'b00001010001100: Data_out <= 16'h1FAC	;
				14'b00001010001101: Data_out <= 16'h1FB8	;
				14'b00001010001110: Data_out <= 16'h1FC4	;
				14'b00001010001111: Data_out <= 16'h1FD1	;
				14'b00001010010000: Data_out <= 16'h1FDD	;
				14'b00001010010001: Data_out <= 16'h1FE9	;
				14'b00001010010010: Data_out <= 16'h1FF5	;
				14'b00001010010011: Data_out <= 16'h2001	;
				14'b00001010010100: Data_out <= 16'h200D	;
				14'b00001010010101: Data_out <= 16'h201A	;
				14'b00001010010110: Data_out <= 16'h2026	;
				14'b00001010010111: Data_out <= 16'h2032	;
				14'b00001010011000: Data_out <= 16'h203E	;
				14'b00001010011001: Data_out <= 16'h204A	;
				14'b00001010011010: Data_out <= 16'h2056	;
				14'b00001010011011: Data_out <= 16'h2063	;
				14'b00001010011100: Data_out <= 16'h206F	;
				14'b00001010011101: Data_out <= 16'h207B	;
				14'b00001010011110: Data_out <= 16'h2087	;
				14'b00001010011111: Data_out <= 16'h2093	;
				14'b00001010100000: Data_out <= 16'h209F	;
				14'b00001010100001: Data_out <= 16'h20AB	;
				14'b00001010100010: Data_out <= 16'h20B8	;
				14'b00001010100011: Data_out <= 16'h20C4	;
				14'b00001010100100: Data_out <= 16'h20D0	;
				14'b00001010100101: Data_out <= 16'h20DC	;
				14'b00001010100110: Data_out <= 16'h20E8	;
				14'b00001010100111: Data_out <= 16'h20F4	;
				14'b00001010101000: Data_out <= 16'h2100	;
				14'b00001010101001: Data_out <= 16'h210D	;
				14'b00001010101010: Data_out <= 16'h2119	;
				14'b00001010101011: Data_out <= 16'h2125	;
				14'b00001010101100: Data_out <= 16'h2131	;
				14'b00001010101101: Data_out <= 16'h213D	;
				14'b00001010101110: Data_out <= 16'h2149	;
				14'b00001010101111: Data_out <= 16'h2155	;
				14'b00001010110000: Data_out <= 16'h2162	;
				14'b00001010110001: Data_out <= 16'h216E	;
				14'b00001010110010: Data_out <= 16'h217A	;
				14'b00001010110011: Data_out <= 16'h2186	;
				14'b00001010110100: Data_out <= 16'h2192	;
				14'b00001010110101: Data_out <= 16'h219E	;
				14'b00001010110110: Data_out <= 16'h21AA	;
				14'b00001010110111: Data_out <= 16'h21B6	;
				14'b00001010111000: Data_out <= 16'h21C3	;
				14'b00001010111001: Data_out <= 16'h21CF	;
				14'b00001010111010: Data_out <= 16'h21DB	;
				14'b00001010111011: Data_out <= 16'h21E7	;
				14'b00001010111100: Data_out <= 16'h21F3	;
				14'b00001010111101: Data_out <= 16'h21FF	;
				14'b00001010111110: Data_out <= 16'h220B	;
				14'b00001010111111: Data_out <= 16'h2217	;
				14'b00001011000000: Data_out <= 16'h2223	;
				14'b00001011000001: Data_out <= 16'h2230	;
				14'b00001011000010: Data_out <= 16'h223C	;
				14'b00001011000011: Data_out <= 16'h2248	;
				14'b00001011000100: Data_out <= 16'h2254	;
				14'b00001011000101: Data_out <= 16'h2260	;
				14'b00001011000110: Data_out <= 16'h226C	;
				14'b00001011000111: Data_out <= 16'h2278	;
				14'b00001011001000: Data_out <= 16'h2284	;
				14'b00001011001001: Data_out <= 16'h2290	;
				14'b00001011001010: Data_out <= 16'h229D	;
				14'b00001011001011: Data_out <= 16'h22A9	;
				14'b00001011001100: Data_out <= 16'h22B5	;
				14'b00001011001101: Data_out <= 16'h22C1	;
				14'b00001011001110: Data_out <= 16'h22CD	;
				14'b00001011001111: Data_out <= 16'h22D9	;
				14'b00001011010000: Data_out <= 16'h22E5	;
				14'b00001011010001: Data_out <= 16'h22F1	;
				14'b00001011010010: Data_out <= 16'h22FD	;
				14'b00001011010011: Data_out <= 16'h2309	;
				14'b00001011010100: Data_out <= 16'h2315	;
				14'b00001011010101: Data_out <= 16'h2322	;
				14'b00001011010110: Data_out <= 16'h232E	;
				14'b00001011010111: Data_out <= 16'h233A	;
				14'b00001011011000: Data_out <= 16'h2346	;
				14'b00001011011001: Data_out <= 16'h2352	;
				14'b00001011011010: Data_out <= 16'h235E	;
				14'b00001011011011: Data_out <= 16'h236A	;
				14'b00001011011100: Data_out <= 16'h2376	;
				14'b00001011011101: Data_out <= 16'h2382	;
				14'b00001011011110: Data_out <= 16'h238E	;
				14'b00001011011111: Data_out <= 16'h239A	;
				14'b00001011100000: Data_out <= 16'h23A6	;
				14'b00001011100001: Data_out <= 16'h23B2	;
				14'b00001011100010: Data_out <= 16'h23BE	;
				14'b00001011100011: Data_out <= 16'h23CB	;
				14'b00001011100100: Data_out <= 16'h23D7	;
				14'b00001011100101: Data_out <= 16'h23E3	;
				14'b00001011100110: Data_out <= 16'h23EF	;
				14'b00001011100111: Data_out <= 16'h23FB	;
				14'b00001011101000: Data_out <= 16'h2407	;
				14'b00001011101001: Data_out <= 16'h2413	;
				14'b00001011101010: Data_out <= 16'h241F	;
				14'b00001011101011: Data_out <= 16'h242B	;
				14'b00001011101100: Data_out <= 16'h2437	;
				14'b00001011101101: Data_out <= 16'h2443	;
				14'b00001011101110: Data_out <= 16'h244F	;
				14'b00001011101111: Data_out <= 16'h245B	;
				14'b00001011110000: Data_out <= 16'h2467	;
				14'b00001011110001: Data_out <= 16'h2473	;
				14'b00001011110010: Data_out <= 16'h247F	;
				14'b00001011110011: Data_out <= 16'h248B	;
				14'b00001011110100: Data_out <= 16'h2497	;
				14'b00001011110101: Data_out <= 16'h24A3	;
				14'b00001011110110: Data_out <= 16'h24B0	;
				14'b00001011110111: Data_out <= 16'h24BC	;
				14'b00001011111000: Data_out <= 16'h24C8	;
				14'b00001011111001: Data_out <= 16'h24D4	;
				14'b00001011111010: Data_out <= 16'h24E0	;
				14'b00001011111011: Data_out <= 16'h24EC	;
				14'b00001011111100: Data_out <= 16'h24F8	;
				14'b00001011111101: Data_out <= 16'h2504	;
				14'b00001011111110: Data_out <= 16'h2510	;
				14'b00001011111111: Data_out <= 16'h251C	;
				14'b00001100000000: Data_out <= 16'h2528	;
				14'b00001100000001: Data_out <= 16'h2534	;
				14'b00001100000010: Data_out <= 16'h2540	;
				14'b00001100000011: Data_out <= 16'h254C	;
				14'b00001100000100: Data_out <= 16'h2558	;
				14'b00001100000101: Data_out <= 16'h2564	;
				14'b00001100000110: Data_out <= 16'h2570	;
				14'b00001100000111: Data_out <= 16'h257C	;
				14'b00001100001000: Data_out <= 16'h2588	;
				14'b00001100001001: Data_out <= 16'h2594	;
				14'b00001100001010: Data_out <= 16'h25A0	;
				14'b00001100001011: Data_out <= 16'h25AC	;
				14'b00001100001100: Data_out <= 16'h25B8	;
				14'b00001100001101: Data_out <= 16'h25C4	;
				14'b00001100001110: Data_out <= 16'h25D0	;
				14'b00001100001111: Data_out <= 16'h25DC	;
				14'b00001100010000: Data_out <= 16'h25E8	;
				14'b00001100010001: Data_out <= 16'h25F4	;
				14'b00001100010010: Data_out <= 16'h2600	;
				14'b00001100010011: Data_out <= 16'h260C	;
				14'b00001100010100: Data_out <= 16'h2618	;
				14'b00001100010101: Data_out <= 16'h2624	;
				14'b00001100010110: Data_out <= 16'h2630	;
				14'b00001100010111: Data_out <= 16'h263C	;
				14'b00001100011000: Data_out <= 16'h2648	;
				14'b00001100011001: Data_out <= 16'h2654	;
				14'b00001100011010: Data_out <= 16'h2660	;
				14'b00001100011011: Data_out <= 16'h266C	;
				14'b00001100011100: Data_out <= 16'h2678	;
				14'b00001100011101: Data_out <= 16'h2684	;
				14'b00001100011110: Data_out <= 16'h2690	;
				14'b00001100011111: Data_out <= 16'h269C	;
				14'b00001100100000: Data_out <= 16'h26A8	;
				14'b00001100100001: Data_out <= 16'h26B4	;
				14'b00001100100010: Data_out <= 16'h26C0	;
				14'b00001100100011: Data_out <= 16'h26CC	;
				14'b00001100100100: Data_out <= 16'h26D8	;
				14'b00001100100101: Data_out <= 16'h26E4	;
				14'b00001100100110: Data_out <= 16'h26F0	;
				14'b00001100100111: Data_out <= 16'h26FC	;
				14'b00001100101000: Data_out <= 16'h2708	;
				14'b00001100101001: Data_out <= 16'h2714	;
				14'b00001100101010: Data_out <= 16'h2720	;
				14'b00001100101011: Data_out <= 16'h272C	;
				14'b00001100101100: Data_out <= 16'h2738	;
				14'b00001100101101: Data_out <= 16'h2744	;
				14'b00001100101110: Data_out <= 16'h274F	;
				14'b00001100101111: Data_out <= 16'h275B	;
				14'b00001100110000: Data_out <= 16'h2767	;
				14'b00001100110001: Data_out <= 16'h2773	;
				14'b00001100110010: Data_out <= 16'h277F	;
				14'b00001100110011: Data_out <= 16'h278B	;
				14'b00001100110100: Data_out <= 16'h2797	;
				14'b00001100110101: Data_out <= 16'h27A3	;
				14'b00001100110110: Data_out <= 16'h27AF	;
				14'b00001100110111: Data_out <= 16'h27BB	;
				14'b00001100111000: Data_out <= 16'h27C7	;
				14'b00001100111001: Data_out <= 16'h27D3	;
				14'b00001100111010: Data_out <= 16'h27DF	;
				14'b00001100111011: Data_out <= 16'h27EB	;
				14'b00001100111100: Data_out <= 16'h27F7	;
				14'b00001100111101: Data_out <= 16'h2803	;
				14'b00001100111110: Data_out <= 16'h280F	;
				14'b00001100111111: Data_out <= 16'h281B	;
				14'b00001101000000: Data_out <= 16'h2827	;
				14'b00001101000001: Data_out <= 16'h2832	;
				14'b00001101000010: Data_out <= 16'h283E	;
				14'b00001101000011: Data_out <= 16'h284A	;
				14'b00001101000100: Data_out <= 16'h2856	;
				14'b00001101000101: Data_out <= 16'h2862	;
				14'b00001101000110: Data_out <= 16'h286E	;
				14'b00001101000111: Data_out <= 16'h287A	;
				14'b00001101001000: Data_out <= 16'h2886	;
				14'b00001101001001: Data_out <= 16'h2892	;
				14'b00001101001010: Data_out <= 16'h289E	;
				14'b00001101001011: Data_out <= 16'h28AA	;
				14'b00001101001100: Data_out <= 16'h28B6	;
				14'b00001101001101: Data_out <= 16'h28C1	;
				14'b00001101001110: Data_out <= 16'h28CD	;
				14'b00001101001111: Data_out <= 16'h28D9	;
				14'b00001101010000: Data_out <= 16'h28E5	;
				14'b00001101010001: Data_out <= 16'h28F1	;
				14'b00001101010010: Data_out <= 16'h28FD	;
				14'b00001101010011: Data_out <= 16'h2909	;
				14'b00001101010100: Data_out <= 16'h2915	;
				14'b00001101010101: Data_out <= 16'h2921	;
				14'b00001101010110: Data_out <= 16'h292D	;
				14'b00001101010111: Data_out <= 16'h2939	;
				14'b00001101011000: Data_out <= 16'h2944	;
				14'b00001101011001: Data_out <= 16'h2950	;
				14'b00001101011010: Data_out <= 16'h295C	;
				14'b00001101011011: Data_out <= 16'h2968	;
				14'b00001101011100: Data_out <= 16'h2974	;
				14'b00001101011101: Data_out <= 16'h2980	;
				14'b00001101011110: Data_out <= 16'h298C	;
				14'b00001101011111: Data_out <= 16'h2998	;
				14'b00001101100000: Data_out <= 16'h29A4	;
				14'b00001101100001: Data_out <= 16'h29AF	;
				14'b00001101100010: Data_out <= 16'h29BB	;
				14'b00001101100011: Data_out <= 16'h29C7	;
				14'b00001101100100: Data_out <= 16'h29D3	;
				14'b00001101100101: Data_out <= 16'h29DF	;
				14'b00001101100110: Data_out <= 16'h29EB	;
				14'b00001101100111: Data_out <= 16'h29F7	;
				14'b00001101101000: Data_out <= 16'h2A03	;
				14'b00001101101001: Data_out <= 16'h2A0E	;
				14'b00001101101010: Data_out <= 16'h2A1A	;
				14'b00001101101011: Data_out <= 16'h2A26	;
				14'b00001101101100: Data_out <= 16'h2A32	;
				14'b00001101101101: Data_out <= 16'h2A3E	;
				14'b00001101101110: Data_out <= 16'h2A4A	;
				14'b00001101101111: Data_out <= 16'h2A56	;
				14'b00001101110000: Data_out <= 16'h2A61	;
				14'b00001101110001: Data_out <= 16'h2A6D	;
				14'b00001101110010: Data_out <= 16'h2A79	;
				14'b00001101110011: Data_out <= 16'h2A85	;
				14'b00001101110100: Data_out <= 16'h2A91	;
				14'b00001101110101: Data_out <= 16'h2A9D	;
				14'b00001101110110: Data_out <= 16'h2AA9	;
				14'b00001101110111: Data_out <= 16'h2AB4	;
				14'b00001101111000: Data_out <= 16'h2AC0	;
				14'b00001101111001: Data_out <= 16'h2ACC	;
				14'b00001101111010: Data_out <= 16'h2AD8	;
				14'b00001101111011: Data_out <= 16'h2AE4	;
				14'b00001101111100: Data_out <= 16'h2AF0	;
				14'b00001101111101: Data_out <= 16'h2AFB	;
				14'b00001101111110: Data_out <= 16'h2B07	;
				14'b00001101111111: Data_out <= 16'h2B13	;
				14'b00001110000000: Data_out <= 16'h2B1F	;
				14'b00001110000001: Data_out <= 16'h2B2B	;
				14'b00001110000010: Data_out <= 16'h2B37	;
				14'b00001110000011: Data_out <= 16'h2B42	;
				14'b00001110000100: Data_out <= 16'h2B4E	;
				14'b00001110000101: Data_out <= 16'h2B5A	;
				14'b00001110000110: Data_out <= 16'h2B66	;
				14'b00001110000111: Data_out <= 16'h2B72	;
				14'b00001110001000: Data_out <= 16'h2B7E	;
				14'b00001110001001: Data_out <= 16'h2B89	;
				14'b00001110001010: Data_out <= 16'h2B95	;
				14'b00001110001011: Data_out <= 16'h2BA1	;
				14'b00001110001100: Data_out <= 16'h2BAD	;
				14'b00001110001101: Data_out <= 16'h2BB9	;
				14'b00001110001110: Data_out <= 16'h2BC4	;
				14'b00001110001111: Data_out <= 16'h2BD0	;
				14'b00001110010000: Data_out <= 16'h2BDC	;
				14'b00001110010001: Data_out <= 16'h2BE8	;
				14'b00001110010010: Data_out <= 16'h2BF4	;
				14'b00001110010011: Data_out <= 16'h2BFF	;
				14'b00001110010100: Data_out <= 16'h2C0B	;
				14'b00001110010101: Data_out <= 16'h2C17	;
				14'b00001110010110: Data_out <= 16'h2C23	;
				14'b00001110010111: Data_out <= 16'h2C2F	;
				14'b00001110011000: Data_out <= 16'h2C3A	;
				14'b00001110011001: Data_out <= 16'h2C46	;
				14'b00001110011010: Data_out <= 16'h2C52	;
				14'b00001110011011: Data_out <= 16'h2C5E	;
				14'b00001110011100: Data_out <= 16'h2C6A	;
				14'b00001110011101: Data_out <= 16'h2C75	;
				14'b00001110011110: Data_out <= 16'h2C81	;
				14'b00001110011111: Data_out <= 16'h2C8D	;
				14'b00001110100000: Data_out <= 16'h2C99	;
				14'b00001110100001: Data_out <= 16'h2CA5	;
				14'b00001110100010: Data_out <= 16'h2CB0	;
				14'b00001110100011: Data_out <= 16'h2CBC	;
				14'b00001110100100: Data_out <= 16'h2CC8	;
				14'b00001110100101: Data_out <= 16'h2CD4	;
				14'b00001110100110: Data_out <= 16'h2CDF	;
				14'b00001110100111: Data_out <= 16'h2CEB	;
				14'b00001110101000: Data_out <= 16'h2CF7	;
				14'b00001110101001: Data_out <= 16'h2D03	;
				14'b00001110101010: Data_out <= 16'h2D0E	;
				14'b00001110101011: Data_out <= 16'h2D1A	;
				14'b00001110101100: Data_out <= 16'h2D26	;
				14'b00001110101101: Data_out <= 16'h2D32	;
				14'b00001110101110: Data_out <= 16'h2D3D	;
				14'b00001110101111: Data_out <= 16'h2D49	;
				14'b00001110110000: Data_out <= 16'h2D55	;
				14'b00001110110001: Data_out <= 16'h2D61	;
				14'b00001110110010: Data_out <= 16'h2D6C	;
				14'b00001110110011: Data_out <= 16'h2D78	;
				14'b00001110110100: Data_out <= 16'h2D84	;
				14'b00001110110101: Data_out <= 16'h2D90	;
				14'b00001110110110: Data_out <= 16'h2D9B	;
				14'b00001110110111: Data_out <= 16'h2DA7	;
				14'b00001110111000: Data_out <= 16'h2DB3	;
				14'b00001110111001: Data_out <= 16'h2DBF	;
				14'b00001110111010: Data_out <= 16'h2DCA	;
				14'b00001110111011: Data_out <= 16'h2DD6	;
				14'b00001110111100: Data_out <= 16'h2DE2	;
				14'b00001110111101: Data_out <= 16'h2DEE	;
				14'b00001110111110: Data_out <= 16'h2DF9	;
				14'b00001110111111: Data_out <= 16'h2E05	;
				14'b00001111000000: Data_out <= 16'h2E11	;
				14'b00001111000001: Data_out <= 16'h2E1D	;
				14'b00001111000010: Data_out <= 16'h2E28	;
				14'b00001111000011: Data_out <= 16'h2E34	;
				14'b00001111000100: Data_out <= 16'h2E40	;
				14'b00001111000101: Data_out <= 16'h2E4B	;
				14'b00001111000110: Data_out <= 16'h2E57	;
				14'b00001111000111: Data_out <= 16'h2E63	;
				14'b00001111001000: Data_out <= 16'h2E6F	;
				14'b00001111001001: Data_out <= 16'h2E7A	;
				14'b00001111001010: Data_out <= 16'h2E86	;
				14'b00001111001011: Data_out <= 16'h2E92	;
				14'b00001111001100: Data_out <= 16'h2E9D	;
				14'b00001111001101: Data_out <= 16'h2EA9	;
				14'b00001111001110: Data_out <= 16'h2EB5	;
				14'b00001111001111: Data_out <= 16'h2EC0	;
				14'b00001111010000: Data_out <= 16'h2ECC	;
				14'b00001111010001: Data_out <= 16'h2ED8	;
				14'b00001111010010: Data_out <= 16'h2EE4	;
				14'b00001111010011: Data_out <= 16'h2EEF	;
				14'b00001111010100: Data_out <= 16'h2EFB	;
				14'b00001111010101: Data_out <= 16'h2F07	;
				14'b00001111010110: Data_out <= 16'h2F12	;
				14'b00001111010111: Data_out <= 16'h2F1E	;
				14'b00001111011000: Data_out <= 16'h2F2A	;
				14'b00001111011001: Data_out <= 16'h2F35	;
				14'b00001111011010: Data_out <= 16'h2F41	;
				14'b00001111011011: Data_out <= 16'h2F4D	;
				14'b00001111011100: Data_out <= 16'h2F58	;
				14'b00001111011101: Data_out <= 16'h2F64	;
				14'b00001111011110: Data_out <= 16'h2F70	;
				14'b00001111011111: Data_out <= 16'h2F7B	;
				14'b00001111100000: Data_out <= 16'h2F87	;
				14'b00001111100001: Data_out <= 16'h2F93	;
				14'b00001111100010: Data_out <= 16'h2F9E	;
				14'b00001111100011: Data_out <= 16'h2FAA	;
				14'b00001111100100: Data_out <= 16'h2FB6	;
				14'b00001111100101: Data_out <= 16'h2FC1	;
				14'b00001111100110: Data_out <= 16'h2FCD	;
				14'b00001111100111: Data_out <= 16'h2FD9	;
				14'b00001111101000: Data_out <= 16'h2FE4	;
				14'b00001111101001: Data_out <= 16'h2FF0	;
				14'b00001111101010: Data_out <= 16'h2FFC	;
				14'b00001111101011: Data_out <= 16'h3007	;
				14'b00001111101100: Data_out <= 16'h3013	;
				14'b00001111101101: Data_out <= 16'h301F	;
				14'b00001111101110: Data_out <= 16'h302A	;
				14'b00001111101111: Data_out <= 16'h3036	;
				14'b00001111110000: Data_out <= 16'h3042	;
				14'b00001111110001: Data_out <= 16'h304D	;
				14'b00001111110010: Data_out <= 16'h3059	;
				14'b00001111110011: Data_out <= 16'h3064	;
				14'b00001111110100: Data_out <= 16'h3070	;
				14'b00001111110101: Data_out <= 16'h307C	;
				14'b00001111110110: Data_out <= 16'h3087	;
				14'b00001111110111: Data_out <= 16'h3093	;
				14'b00001111111000: Data_out <= 16'h309F	;
				14'b00001111111001: Data_out <= 16'h30AA	;
				14'b00001111111010: Data_out <= 16'h30B6	;
				14'b00001111111011: Data_out <= 16'h30C1	;
				14'b00001111111100: Data_out <= 16'h30CD	;
				14'b00001111111101: Data_out <= 16'h30D9	;
				14'b00001111111110: Data_out <= 16'h30E4	;
				14'b00001111111111: Data_out <= 16'h30F0	;
				14'b00010000000000: Data_out <= 16'h30FB	;
				14'b00010000000001: Data_out <= 16'h3107	;
				14'b00010000000010: Data_out <= 16'h3113	;
				14'b00010000000011: Data_out <= 16'h311E	;
				14'b00010000000100: Data_out <= 16'h312A	;
				14'b00010000000101: Data_out <= 16'h3136	;
				14'b00010000000110: Data_out <= 16'h3141	;
				14'b00010000000111: Data_out <= 16'h314D	;
				14'b00010000001000: Data_out <= 16'h3158	;
				14'b00010000001001: Data_out <= 16'h3164	;
				14'b00010000001010: Data_out <= 16'h316F	;
				14'b00010000001011: Data_out <= 16'h317B	;
				14'b00010000001100: Data_out <= 16'h3187	;
				14'b00010000001101: Data_out <= 16'h3192	;
				14'b00010000001110: Data_out <= 16'h319E	;
				14'b00010000001111: Data_out <= 16'h31A9	;
				14'b00010000010000: Data_out <= 16'h31B5	;
				14'b00010000010001: Data_out <= 16'h31C1	;
				14'b00010000010010: Data_out <= 16'h31CC	;
				14'b00010000010011: Data_out <= 16'h31D8	;
				14'b00010000010100: Data_out <= 16'h31E3	;
				14'b00010000010101: Data_out <= 16'h31EF	;
				14'b00010000010110: Data_out <= 16'h31FA	;
				14'b00010000010111: Data_out <= 16'h3206	;
				14'b00010000011000: Data_out <= 16'h3212	;
				14'b00010000011001: Data_out <= 16'h321D	;
				14'b00010000011010: Data_out <= 16'h3229	;
				14'b00010000011011: Data_out <= 16'h3234	;
				14'b00010000011100: Data_out <= 16'h3240	;
				14'b00010000011101: Data_out <= 16'h324B	;
				14'b00010000011110: Data_out <= 16'h3257	;
				14'b00010000011111: Data_out <= 16'h3262	;
				14'b00010000100000: Data_out <= 16'h326E	;
				14'b00010000100001: Data_out <= 16'h327A	;
				14'b00010000100010: Data_out <= 16'h3285	;
				14'b00010000100011: Data_out <= 16'h3291	;
				14'b00010000100100: Data_out <= 16'h329C	;
				14'b00010000100101: Data_out <= 16'h32A8	;
				14'b00010000100110: Data_out <= 16'h32B3	;
				14'b00010000100111: Data_out <= 16'h32BF	;
				14'b00010000101000: Data_out <= 16'h32CA	;
				14'b00010000101001: Data_out <= 16'h32D6	;
				14'b00010000101010: Data_out <= 16'h32E1	;
				14'b00010000101011: Data_out <= 16'h32ED	;
				14'b00010000101100: Data_out <= 16'h32F8	;
				14'b00010000101101: Data_out <= 16'h3304	;
				14'b00010000101110: Data_out <= 16'h3310	;
				14'b00010000101111: Data_out <= 16'h331B	;
				14'b00010000110000: Data_out <= 16'h3327	;
				14'b00010000110001: Data_out <= 16'h3332	;
				14'b00010000110010: Data_out <= 16'h333E	;
				14'b00010000110011: Data_out <= 16'h3349	;
				14'b00010000110100: Data_out <= 16'h3355	;
				14'b00010000110101: Data_out <= 16'h3360	;
				14'b00010000110110: Data_out <= 16'h336C	;
				14'b00010000110111: Data_out <= 16'h3377	;
				14'b00010000111000: Data_out <= 16'h3383	;
				14'b00010000111001: Data_out <= 16'h338E	;
				14'b00010000111010: Data_out <= 16'h339A	;
				14'b00010000111011: Data_out <= 16'h33A5	;
				14'b00010000111100: Data_out <= 16'h33B1	;
				14'b00010000111101: Data_out <= 16'h33BC	;
				14'b00010000111110: Data_out <= 16'h33C8	;
				14'b00010000111111: Data_out <= 16'h33D3	;
				14'b00010001000000: Data_out <= 16'h33DF	;
				14'b00010001000001: Data_out <= 16'h33EA	;
				14'b00010001000010: Data_out <= 16'h33F6	;
				14'b00010001000011: Data_out <= 16'h3401	;
				14'b00010001000100: Data_out <= 16'h340D	;
				14'b00010001000101: Data_out <= 16'h3418	;
				14'b00010001000110: Data_out <= 16'h3424	;
				14'b00010001000111: Data_out <= 16'h342F	;
				14'b00010001001000: Data_out <= 16'h343A	;
				14'b00010001001001: Data_out <= 16'h3446	;
				14'b00010001001010: Data_out <= 16'h3451	;
				14'b00010001001011: Data_out <= 16'h345D	;
				14'b00010001001100: Data_out <= 16'h3468	;
				14'b00010001001101: Data_out <= 16'h3474	;
				14'b00010001001110: Data_out <= 16'h347F	;
				14'b00010001001111: Data_out <= 16'h348B	;
				14'b00010001010000: Data_out <= 16'h3496	;
				14'b00010001010001: Data_out <= 16'h34A2	;
				14'b00010001010010: Data_out <= 16'h34AD	;
				14'b00010001010011: Data_out <= 16'h34B9	;
				14'b00010001010100: Data_out <= 16'h34C4	;
				14'b00010001010101: Data_out <= 16'h34CF	;
				14'b00010001010110: Data_out <= 16'h34DB	;
				14'b00010001010111: Data_out <= 16'h34E6	;
				14'b00010001011000: Data_out <= 16'h34F2	;
				14'b00010001011001: Data_out <= 16'h34FD	;
				14'b00010001011010: Data_out <= 16'h3509	;
				14'b00010001011011: Data_out <= 16'h3514	;
				14'b00010001011100: Data_out <= 16'h3520	;
				14'b00010001011101: Data_out <= 16'h352B	;
				14'b00010001011110: Data_out <= 16'h3536	;
				14'b00010001011111: Data_out <= 16'h3542	;
				14'b00010001100000: Data_out <= 16'h354D	;
				14'b00010001100001: Data_out <= 16'h3559	;
				14'b00010001100010: Data_out <= 16'h3564	;
				14'b00010001100011: Data_out <= 16'h3570	;
				14'b00010001100100: Data_out <= 16'h357B	;
				14'b00010001100101: Data_out <= 16'h3586	;
				14'b00010001100110: Data_out <= 16'h3592	;
				14'b00010001100111: Data_out <= 16'h359D	;
				14'b00010001101000: Data_out <= 16'h35A9	;
				14'b00010001101001: Data_out <= 16'h35B4	;
				14'b00010001101010: Data_out <= 16'h35BF	;
				14'b00010001101011: Data_out <= 16'h35CB	;
				14'b00010001101100: Data_out <= 16'h35D6	;
				14'b00010001101101: Data_out <= 16'h35E2	;
				14'b00010001101110: Data_out <= 16'h35ED	;
				14'b00010001101111: Data_out <= 16'h35F8	;
				14'b00010001110000: Data_out <= 16'h3604	;
				14'b00010001110001: Data_out <= 16'h360F	;
				14'b00010001110010: Data_out <= 16'h361B	;
				14'b00010001110011: Data_out <= 16'h3626	;
				14'b00010001110100: Data_out <= 16'h3631	;
				14'b00010001110101: Data_out <= 16'h363D	;
				14'b00010001110110: Data_out <= 16'h3648	;
				14'b00010001110111: Data_out <= 16'h3653	;
				14'b00010001111000: Data_out <= 16'h365F	;
				14'b00010001111001: Data_out <= 16'h366A	;
				14'b00010001111010: Data_out <= 16'h3676	;
				14'b00010001111011: Data_out <= 16'h3681	;
				14'b00010001111100: Data_out <= 16'h368C	;
				14'b00010001111101: Data_out <= 16'h3698	;
				14'b00010001111110: Data_out <= 16'h36A3	;
				14'b00010001111111: Data_out <= 16'h36AE	;
				14'b00010010000000: Data_out <= 16'h36BA	;
				14'b00010010000001: Data_out <= 16'h36C5	;
				14'b00010010000010: Data_out <= 16'h36D1	;
				14'b00010010000011: Data_out <= 16'h36DC	;
				14'b00010010000100: Data_out <= 16'h36E7	;
				14'b00010010000101: Data_out <= 16'h36F3	;
				14'b00010010000110: Data_out <= 16'h36FE	;
				14'b00010010000111: Data_out <= 16'h3709	;
				14'b00010010001000: Data_out <= 16'h3715	;
				14'b00010010001001: Data_out <= 16'h3720	;
				14'b00010010001010: Data_out <= 16'h372B	;
				14'b00010010001011: Data_out <= 16'h3737	;
				14'b00010010001100: Data_out <= 16'h3742	;
				14'b00010010001101: Data_out <= 16'h374D	;
				14'b00010010001110: Data_out <= 16'h3759	;
				14'b00010010001111: Data_out <= 16'h3764	;
				14'b00010010010000: Data_out <= 16'h376F	;
				14'b00010010010001: Data_out <= 16'h377B	;
				14'b00010010010010: Data_out <= 16'h3786	;
				14'b00010010010011: Data_out <= 16'h3791	;
				14'b00010010010100: Data_out <= 16'h379D	;
				14'b00010010010101: Data_out <= 16'h37A8	;
				14'b00010010010110: Data_out <= 16'h37B3	;
				14'b00010010010111: Data_out <= 16'h37BF	;
				14'b00010010011000: Data_out <= 16'h37CA	;
				14'b00010010011001: Data_out <= 16'h37D5	;
				14'b00010010011010: Data_out <= 16'h37E0	;
				14'b00010010011011: Data_out <= 16'h37EC	;
				14'b00010010011100: Data_out <= 16'h37F7	;
				14'b00010010011101: Data_out <= 16'h3802	;
				14'b00010010011110: Data_out <= 16'h380E	;
				14'b00010010011111: Data_out <= 16'h3819	;
				14'b00010010100000: Data_out <= 16'h3824	;
				14'b00010010100001: Data_out <= 16'h3830	;
				14'b00010010100010: Data_out <= 16'h383B	;
				14'b00010010100011: Data_out <= 16'h3846	;
				14'b00010010100100: Data_out <= 16'h3851	;
				14'b00010010100101: Data_out <= 16'h385D	;
				14'b00010010100110: Data_out <= 16'h3868	;
				14'b00010010100111: Data_out <= 16'h3873	;
				14'b00010010101000: Data_out <= 16'h387F	;
				14'b00010010101001: Data_out <= 16'h388A	;
				14'b00010010101010: Data_out <= 16'h3895	;
				14'b00010010101011: Data_out <= 16'h38A0	;
				14'b00010010101100: Data_out <= 16'h38AC	;
				14'b00010010101101: Data_out <= 16'h38B7	;
				14'b00010010101110: Data_out <= 16'h38C2	;
				14'b00010010101111: Data_out <= 16'h38CD	;
				14'b00010010110000: Data_out <= 16'h38D9	;
				14'b00010010110001: Data_out <= 16'h38E4	;
				14'b00010010110010: Data_out <= 16'h38EF	;
				14'b00010010110011: Data_out <= 16'h38FA	;
				14'b00010010110100: Data_out <= 16'h3906	;
				14'b00010010110101: Data_out <= 16'h3911	;
				14'b00010010110110: Data_out <= 16'h391C	;
				14'b00010010110111: Data_out <= 16'h3927	;
				14'b00010010111000: Data_out <= 16'h3933	;
				14'b00010010111001: Data_out <= 16'h393E	;
				14'b00010010111010: Data_out <= 16'h3949	;
				14'b00010010111011: Data_out <= 16'h3954	;
				14'b00010010111100: Data_out <= 16'h3960	;
				14'b00010010111101: Data_out <= 16'h396B	;
				14'b00010010111110: Data_out <= 16'h3976	;
				14'b00010010111111: Data_out <= 16'h3981	;
				14'b00010011000000: Data_out <= 16'h398D	;
				14'b00010011000001: Data_out <= 16'h3998	;
				14'b00010011000010: Data_out <= 16'h39A3	;
				14'b00010011000011: Data_out <= 16'h39AE	;
				14'b00010011000100: Data_out <= 16'h39B9	;
				14'b00010011000101: Data_out <= 16'h39C5	;
				14'b00010011000110: Data_out <= 16'h39D0	;
				14'b00010011000111: Data_out <= 16'h39DB	;
				14'b00010011001000: Data_out <= 16'h39E6	;
				14'b00010011001001: Data_out <= 16'h39F1	;
				14'b00010011001010: Data_out <= 16'h39FD	;
				14'b00010011001011: Data_out <= 16'h3A08	;
				14'b00010011001100: Data_out <= 16'h3A13	;
				14'b00010011001101: Data_out <= 16'h3A1E	;
				14'b00010011001110: Data_out <= 16'h3A29	;
				14'b00010011001111: Data_out <= 16'h3A35	;
				14'b00010011010000: Data_out <= 16'h3A40	;
				14'b00010011010001: Data_out <= 16'h3A4B	;
				14'b00010011010010: Data_out <= 16'h3A56	;
				14'b00010011010011: Data_out <= 16'h3A61	;
				14'b00010011010100: Data_out <= 16'h3A6D	;
				14'b00010011010101: Data_out <= 16'h3A78	;
				14'b00010011010110: Data_out <= 16'h3A83	;
				14'b00010011010111: Data_out <= 16'h3A8E	;
				14'b00010011011000: Data_out <= 16'h3A99	;
				14'b00010011011001: Data_out <= 16'h3AA4	;
				14'b00010011011010: Data_out <= 16'h3AB0	;
				14'b00010011011011: Data_out <= 16'h3ABB	;
				14'b00010011011100: Data_out <= 16'h3AC6	;
				14'b00010011011101: Data_out <= 16'h3AD1	;
				14'b00010011011110: Data_out <= 16'h3ADC	;
				14'b00010011011111: Data_out <= 16'h3AE7	;
				14'b00010011100000: Data_out <= 16'h3AF3	;
				14'b00010011100001: Data_out <= 16'h3AFE	;
				14'b00010011100010: Data_out <= 16'h3B09	;
				14'b00010011100011: Data_out <= 16'h3B14	;
				14'b00010011100100: Data_out <= 16'h3B1F	;
				14'b00010011100101: Data_out <= 16'h3B2A	;
				14'b00010011100110: Data_out <= 16'h3B35	;
				14'b00010011100111: Data_out <= 16'h3B41	;
				14'b00010011101000: Data_out <= 16'h3B4C	;
				14'b00010011101001: Data_out <= 16'h3B57	;
				14'b00010011101010: Data_out <= 16'h3B62	;
				14'b00010011101011: Data_out <= 16'h3B6D	;
				14'b00010011101100: Data_out <= 16'h3B78	;
				14'b00010011101101: Data_out <= 16'h3B83	;
				14'b00010011101110: Data_out <= 16'h3B8F	;
				14'b00010011101111: Data_out <= 16'h3B9A	;
				14'b00010011110000: Data_out <= 16'h3BA5	;
				14'b00010011110001: Data_out <= 16'h3BB0	;
				14'b00010011110010: Data_out <= 16'h3BBB	;
				14'b00010011110011: Data_out <= 16'h3BC6	;
				14'b00010011110100: Data_out <= 16'h3BD1	;
				14'b00010011110101: Data_out <= 16'h3BDC	;
				14'b00010011110110: Data_out <= 16'h3BE7	;
				14'b00010011110111: Data_out <= 16'h3BF3	;
				14'b00010011111000: Data_out <= 16'h3BFE	;
				14'b00010011111001: Data_out <= 16'h3C09	;
				14'b00010011111010: Data_out <= 16'h3C14	;
				14'b00010011111011: Data_out <= 16'h3C1F	;
				14'b00010011111100: Data_out <= 16'h3C2A	;
				14'b00010011111101: Data_out <= 16'h3C35	;
				14'b00010011111110: Data_out <= 16'h3C40	;
				14'b00010011111111: Data_out <= 16'h3C4B	;
				14'b00010100000000: Data_out <= 16'h3C56	;
				14'b00010100000001: Data_out <= 16'h3C61	;
				14'b00010100000010: Data_out <= 16'h3C6D	;
				14'b00010100000011: Data_out <= 16'h3C78	;
				14'b00010100000100: Data_out <= 16'h3C83	;
				14'b00010100000101: Data_out <= 16'h3C8E	;
				14'b00010100000110: Data_out <= 16'h3C99	;
				14'b00010100000111: Data_out <= 16'h3CA4	;
				14'b00010100001000: Data_out <= 16'h3CAF	;
				14'b00010100001001: Data_out <= 16'h3CBA	;
				14'b00010100001010: Data_out <= 16'h3CC5	;
				14'b00010100001011: Data_out <= 16'h3CD0	;
				14'b00010100001100: Data_out <= 16'h3CDB	;
				14'b00010100001101: Data_out <= 16'h3CE6	;
				14'b00010100001110: Data_out <= 16'h3CF1	;
				14'b00010100001111: Data_out <= 16'h3CFC	;
				14'b00010100010000: Data_out <= 16'h3D07	;
				14'b00010100010001: Data_out <= 16'h3D12	;
				14'b00010100010010: Data_out <= 16'h3D1D	;
				14'b00010100010011: Data_out <= 16'h3D29	;
				14'b00010100010100: Data_out <= 16'h3D34	;
				14'b00010100010101: Data_out <= 16'h3D3F	;
				14'b00010100010110: Data_out <= 16'h3D4A	;
				14'b00010100010111: Data_out <= 16'h3D55	;
				14'b00010100011000: Data_out <= 16'h3D60	;
				14'b00010100011001: Data_out <= 16'h3D6B	;
				14'b00010100011010: Data_out <= 16'h3D76	;
				14'b00010100011011: Data_out <= 16'h3D81	;
				14'b00010100011100: Data_out <= 16'h3D8C	;
				14'b00010100011101: Data_out <= 16'h3D97	;
				14'b00010100011110: Data_out <= 16'h3DA2	;
				14'b00010100011111: Data_out <= 16'h3DAD	;
				14'b00010100100000: Data_out <= 16'h3DB8	;
				14'b00010100100001: Data_out <= 16'h3DC3	;
				14'b00010100100010: Data_out <= 16'h3DCE	;
				14'b00010100100011: Data_out <= 16'h3DD9	;
				14'b00010100100100: Data_out <= 16'h3DE4	;
				14'b00010100100101: Data_out <= 16'h3DEF	;
				14'b00010100100110: Data_out <= 16'h3DFA	;
				14'b00010100100111: Data_out <= 16'h3E05	;
				14'b00010100101000: Data_out <= 16'h3E10	;
				14'b00010100101001: Data_out <= 16'h3E1B	;
				14'b00010100101010: Data_out <= 16'h3E26	;
				14'b00010100101011: Data_out <= 16'h3E31	;
				14'b00010100101100: Data_out <= 16'h3E3C	;
				14'b00010100101101: Data_out <= 16'h3E47	;
				14'b00010100101110: Data_out <= 16'h3E52	;
				14'b00010100101111: Data_out <= 16'h3E5D	;
				14'b00010100110000: Data_out <= 16'h3E68	;
				14'b00010100110001: Data_out <= 16'h3E73	;
				14'b00010100110010: Data_out <= 16'h3E7E	;
				14'b00010100110011: Data_out <= 16'h3E89	;
				14'b00010100110100: Data_out <= 16'h3E94	;
				14'b00010100110101: Data_out <= 16'h3E9E	;
				14'b00010100110110: Data_out <= 16'h3EA9	;
				14'b00010100110111: Data_out <= 16'h3EB4	;
				14'b00010100111000: Data_out <= 16'h3EBF	;
				14'b00010100111001: Data_out <= 16'h3ECA	;
				14'b00010100111010: Data_out <= 16'h3ED5	;
				14'b00010100111011: Data_out <= 16'h3EE0	;
				14'b00010100111100: Data_out <= 16'h3EEB	;
				14'b00010100111101: Data_out <= 16'h3EF6	;
				14'b00010100111110: Data_out <= 16'h3F01	;
				14'b00010100111111: Data_out <= 16'h3F0C	;
				14'b00010101000000: Data_out <= 16'h3F17	;
				14'b00010101000001: Data_out <= 16'h3F22	;
				14'b00010101000010: Data_out <= 16'h3F2D	;
				14'b00010101000011: Data_out <= 16'h3F38	;
				14'b00010101000100: Data_out <= 16'h3F43	;
				14'b00010101000101: Data_out <= 16'h3F4E	;
				14'b00010101000110: Data_out <= 16'h3F58	;
				14'b00010101000111: Data_out <= 16'h3F63	;
				14'b00010101001000: Data_out <= 16'h3F6E	;
				14'b00010101001001: Data_out <= 16'h3F79	;
				14'b00010101001010: Data_out <= 16'h3F84	;
				14'b00010101001011: Data_out <= 16'h3F8F	;
				14'b00010101001100: Data_out <= 16'h3F9A	;
				14'b00010101001101: Data_out <= 16'h3FA5	;
				14'b00010101001110: Data_out <= 16'h3FB0	;
				14'b00010101001111: Data_out <= 16'h3FBB	;
				14'b00010101010000: Data_out <= 16'h3FC6	;
				14'b00010101010001: Data_out <= 16'h3FD0	;
				14'b00010101010010: Data_out <= 16'h3FDB	;
				14'b00010101010011: Data_out <= 16'h3FE6	;
				14'b00010101010100: Data_out <= 16'h3FF1	;
				14'b00010101010101: Data_out <= 16'h3FFC	;
				14'b00010101010110: Data_out <= 16'h4007	;
				14'b00010101010111: Data_out <= 16'h4012	;
				14'b00010101011000: Data_out <= 16'h401D	;
				14'b00010101011001: Data_out <= 16'h4027	;
				14'b00010101011010: Data_out <= 16'h4032	;
				14'b00010101011011: Data_out <= 16'h403D	;
				14'b00010101011100: Data_out <= 16'h4048	;
				14'b00010101011101: Data_out <= 16'h4053	;
				14'b00010101011110: Data_out <= 16'h405E	;
				14'b00010101011111: Data_out <= 16'h4069	;
				14'b00010101100000: Data_out <= 16'h4074	;
				14'b00010101100001: Data_out <= 16'h407E	;
				14'b00010101100010: Data_out <= 16'h4089	;
				14'b00010101100011: Data_out <= 16'h4094	;
				14'b00010101100100: Data_out <= 16'h409F	;
				14'b00010101100101: Data_out <= 16'h40AA	;
				14'b00010101100110: Data_out <= 16'h40B5	;
				14'b00010101100111: Data_out <= 16'h40BF	;
				14'b00010101101000: Data_out <= 16'h40CA	;
				14'b00010101101001: Data_out <= 16'h40D5	;
				14'b00010101101010: Data_out <= 16'h40E0	;
				14'b00010101101011: Data_out <= 16'h40EB	;
				14'b00010101101100: Data_out <= 16'h40F6	;
				14'b00010101101101: Data_out <= 16'h4100	;
				14'b00010101101110: Data_out <= 16'h410B	;
				14'b00010101101111: Data_out <= 16'h4116	;
				14'b00010101110000: Data_out <= 16'h4121	;
				14'b00010101110001: Data_out <= 16'h412C	;
				14'b00010101110010: Data_out <= 16'h4137	;
				14'b00010101110011: Data_out <= 16'h4141	;
				14'b00010101110100: Data_out <= 16'h414C	;
				14'b00010101110101: Data_out <= 16'h4157	;
				14'b00010101110110: Data_out <= 16'h4162	;
				14'b00010101110111: Data_out <= 16'h416D	;
				14'b00010101111000: Data_out <= 16'h4177	;
				14'b00010101111001: Data_out <= 16'h4182	;
				14'b00010101111010: Data_out <= 16'h418D	;
				14'b00010101111011: Data_out <= 16'h4198	;
				14'b00010101111100: Data_out <= 16'h41A3	;
				14'b00010101111101: Data_out <= 16'h41AD	;
				14'b00010101111110: Data_out <= 16'h41B8	;
				14'b00010101111111: Data_out <= 16'h41C3	;
				14'b00010110000000: Data_out <= 16'h41CE	;
				14'b00010110000001: Data_out <= 16'h41D8	;
				14'b00010110000010: Data_out <= 16'h41E3	;
				14'b00010110000011: Data_out <= 16'h41EE	;
				14'b00010110000100: Data_out <= 16'h41F9	;
				14'b00010110000101: Data_out <= 16'h4204	;
				14'b00010110000110: Data_out <= 16'h420E	;
				14'b00010110000111: Data_out <= 16'h4219	;
				14'b00010110001000: Data_out <= 16'h4224	;
				14'b00010110001001: Data_out <= 16'h422F	;
				14'b00010110001010: Data_out <= 16'h4239	;
				14'b00010110001011: Data_out <= 16'h4244	;
				14'b00010110001100: Data_out <= 16'h424F	;
				14'b00010110001101: Data_out <= 16'h425A	;
				14'b00010110001110: Data_out <= 16'h4264	;
				14'b00010110001111: Data_out <= 16'h426F	;
				14'b00010110010000: Data_out <= 16'h427A	;
				14'b00010110010001: Data_out <= 16'h4285	;
				14'b00010110010010: Data_out <= 16'h428F	;
				14'b00010110010011: Data_out <= 16'h429A	;
				14'b00010110010100: Data_out <= 16'h42A5	;
				14'b00010110010101: Data_out <= 16'h42AF	;
				14'b00010110010110: Data_out <= 16'h42BA	;
				14'b00010110010111: Data_out <= 16'h42C5	;
				14'b00010110011000: Data_out <= 16'h42D0	;
				14'b00010110011001: Data_out <= 16'h42DA	;
				14'b00010110011010: Data_out <= 16'h42E5	;
				14'b00010110011011: Data_out <= 16'h42F0	;
				14'b00010110011100: Data_out <= 16'h42FB	;
				14'b00010110011101: Data_out <= 16'h4305	;
				14'b00010110011110: Data_out <= 16'h4310	;
				14'b00010110011111: Data_out <= 16'h431B	;
				14'b00010110100000: Data_out <= 16'h4325	;
				14'b00010110100001: Data_out <= 16'h4330	;
				14'b00010110100010: Data_out <= 16'h433B	;
				14'b00010110100011: Data_out <= 16'h4345	;
				14'b00010110100100: Data_out <= 16'h4350	;
				14'b00010110100101: Data_out <= 16'h435B	;
				14'b00010110100110: Data_out <= 16'h4365	;
				14'b00010110100111: Data_out <= 16'h4370	;
				14'b00010110101000: Data_out <= 16'h437B	;
				14'b00010110101001: Data_out <= 16'h4386	;
				14'b00010110101010: Data_out <= 16'h4390	;
				14'b00010110101011: Data_out <= 16'h439B	;
				14'b00010110101100: Data_out <= 16'h43A6	;
				14'b00010110101101: Data_out <= 16'h43B0	;
				14'b00010110101110: Data_out <= 16'h43BB	;
				14'b00010110101111: Data_out <= 16'h43C6	;
				14'b00010110110000: Data_out <= 16'h43D0	;
				14'b00010110110001: Data_out <= 16'h43DB	;
				14'b00010110110010: Data_out <= 16'h43E5	;
				14'b00010110110011: Data_out <= 16'h43F0	;
				14'b00010110110100: Data_out <= 16'h43FB	;
				14'b00010110110101: Data_out <= 16'h4405	;
				14'b00010110110110: Data_out <= 16'h4410	;
				14'b00010110110111: Data_out <= 16'h441B	;
				14'b00010110111000: Data_out <= 16'h4425	;
				14'b00010110111001: Data_out <= 16'h4430	;
				14'b00010110111010: Data_out <= 16'h443B	;
				14'b00010110111011: Data_out <= 16'h4445	;
				14'b00010110111100: Data_out <= 16'h4450	;
				14'b00010110111101: Data_out <= 16'h445B	;
				14'b00010110111110: Data_out <= 16'h4465	;
				14'b00010110111111: Data_out <= 16'h4470	;
				14'b00010111000000: Data_out <= 16'h447A	;
				14'b00010111000001: Data_out <= 16'h4485	;
				14'b00010111000010: Data_out <= 16'h4490	;
				14'b00010111000011: Data_out <= 16'h449A	;
				14'b00010111000100: Data_out <= 16'h44A5	;
				14'b00010111000101: Data_out <= 16'h44AF	;
				14'b00010111000110: Data_out <= 16'h44BA	;
				14'b00010111000111: Data_out <= 16'h44C5	;
				14'b00010111001000: Data_out <= 16'h44CF	;
				14'b00010111001001: Data_out <= 16'h44DA	;
				14'b00010111001010: Data_out <= 16'h44E4	;
				14'b00010111001011: Data_out <= 16'h44EF	;
				14'b00010111001100: Data_out <= 16'h44FA	;
				14'b00010111001101: Data_out <= 16'h4504	;
				14'b00010111001110: Data_out <= 16'h450F	;
				14'b00010111001111: Data_out <= 16'h4519	;
				14'b00010111010000: Data_out <= 16'h4524	;
				14'b00010111010001: Data_out <= 16'h452E	;
				14'b00010111010010: Data_out <= 16'h4539	;
				14'b00010111010011: Data_out <= 16'h4544	;
				14'b00010111010100: Data_out <= 16'h454E	;
				14'b00010111010101: Data_out <= 16'h4559	;
				14'b00010111010110: Data_out <= 16'h4563	;
				14'b00010111010111: Data_out <= 16'h456E	;
				14'b00010111011000: Data_out <= 16'h4578	;
				14'b00010111011001: Data_out <= 16'h4583	;
				14'b00010111011010: Data_out <= 16'h458E	;
				14'b00010111011011: Data_out <= 16'h4598	;
				14'b00010111011100: Data_out <= 16'h45A3	;
				14'b00010111011101: Data_out <= 16'h45AD	;
				14'b00010111011110: Data_out <= 16'h45B8	;
				14'b00010111011111: Data_out <= 16'h45C2	;
				14'b00010111100000: Data_out <= 16'h45CD	;
				14'b00010111100001: Data_out <= 16'h45D7	;
				14'b00010111100010: Data_out <= 16'h45E2	;
				14'b00010111100011: Data_out <= 16'h45EC	;
				14'b00010111100100: Data_out <= 16'h45F7	;
				14'b00010111100101: Data_out <= 16'h4601	;
				14'b00010111100110: Data_out <= 16'h460C	;
				14'b00010111100111: Data_out <= 16'h4616	;
				14'b00010111101000: Data_out <= 16'h4621	;
				14'b00010111101001: Data_out <= 16'h462B	;
				14'b00010111101010: Data_out <= 16'h4636	;
				14'b00010111101011: Data_out <= 16'h4640	;
				14'b00010111101100: Data_out <= 16'h464B	;
				14'b00010111101101: Data_out <= 16'h4655	;
				14'b00010111101110: Data_out <= 16'h4660	;
				14'b00010111101111: Data_out <= 16'h466A	;
				14'b00010111110000: Data_out <= 16'h4675	;
				14'b00010111110001: Data_out <= 16'h467F	;
				14'b00010111110010: Data_out <= 16'h468A	;
				14'b00010111110011: Data_out <= 16'h4694	;
				14'b00010111110100: Data_out <= 16'h469F	;
				14'b00010111110101: Data_out <= 16'h46A9	;
				14'b00010111110110: Data_out <= 16'h46B4	;
				14'b00010111110111: Data_out <= 16'h46BE	;
				14'b00010111111000: Data_out <= 16'h46C9	;
				14'b00010111111001: Data_out <= 16'h46D3	;
				14'b00010111111010: Data_out <= 16'h46DE	;
				14'b00010111111011: Data_out <= 16'h46E8	;
				14'b00010111111100: Data_out <= 16'h46F3	;
				14'b00010111111101: Data_out <= 16'h46FD	;
				14'b00010111111110: Data_out <= 16'h4708	;
				14'b00010111111111: Data_out <= 16'h4712	;
				14'b00011000000000: Data_out <= 16'h471C	;
				14'b00011000000001: Data_out <= 16'h4727	;
				14'b00011000000010: Data_out <= 16'h4731	;
				14'b00011000000011: Data_out <= 16'h473C	;
				14'b00011000000100: Data_out <= 16'h4746	;
				14'b00011000000101: Data_out <= 16'h4751	;
				14'b00011000000110: Data_out <= 16'h475B	;
				14'b00011000000111: Data_out <= 16'h4766	;
				14'b00011000001000: Data_out <= 16'h4770	;
				14'b00011000001001: Data_out <= 16'h477A	;
				14'b00011000001010: Data_out <= 16'h4785	;
				14'b00011000001011: Data_out <= 16'h478F	;
				14'b00011000001100: Data_out <= 16'h479A	;
				14'b00011000001101: Data_out <= 16'h47A4	;
				14'b00011000001110: Data_out <= 16'h47AE	;
				14'b00011000001111: Data_out <= 16'h47B9	;
				14'b00011000010000: Data_out <= 16'h47C3	;
				14'b00011000010001: Data_out <= 16'h47CE	;
				14'b00011000010010: Data_out <= 16'h47D8	;
				14'b00011000010011: Data_out <= 16'h47E3	;
				14'b00011000010100: Data_out <= 16'h47ED	;
				14'b00011000010101: Data_out <= 16'h47F7	;
				14'b00011000010110: Data_out <= 16'h4802	;
				14'b00011000010111: Data_out <= 16'h480C	;
				14'b00011000011000: Data_out <= 16'h4816	;
				14'b00011000011001: Data_out <= 16'h4821	;
				14'b00011000011010: Data_out <= 16'h482B	;
				14'b00011000011011: Data_out <= 16'h4836	;
				14'b00011000011100: Data_out <= 16'h4840	;
				14'b00011000011101: Data_out <= 16'h484A	;
				14'b00011000011110: Data_out <= 16'h4855	;
				14'b00011000011111: Data_out <= 16'h485F	;
				14'b00011000100000: Data_out <= 16'h4869	;
				14'b00011000100001: Data_out <= 16'h4874	;
				14'b00011000100010: Data_out <= 16'h487E	;
				14'b00011000100011: Data_out <= 16'h4889	;
				14'b00011000100100: Data_out <= 16'h4893	;
				14'b00011000100101: Data_out <= 16'h489D	;
				14'b00011000100110: Data_out <= 16'h48A8	;
				14'b00011000100111: Data_out <= 16'h48B2	;
				14'b00011000101000: Data_out <= 16'h48BC	;
				14'b00011000101001: Data_out <= 16'h48C7	;
				14'b00011000101010: Data_out <= 16'h48D1	;
				14'b00011000101011: Data_out <= 16'h48DB	;
				14'b00011000101100: Data_out <= 16'h48E6	;
				14'b00011000101101: Data_out <= 16'h48F0	;
				14'b00011000101110: Data_out <= 16'h48FA	;
				14'b00011000101111: Data_out <= 16'h4905	;
				14'b00011000110000: Data_out <= 16'h490F	;
				14'b00011000110001: Data_out <= 16'h4919	;
				14'b00011000110010: Data_out <= 16'h4924	;
				14'b00011000110011: Data_out <= 16'h492E	;
				14'b00011000110100: Data_out <= 16'h4938	;
				14'b00011000110101: Data_out <= 16'h4942	;
				14'b00011000110110: Data_out <= 16'h494D	;
				14'b00011000110111: Data_out <= 16'h4957	;
				14'b00011000111000: Data_out <= 16'h4961	;
				14'b00011000111001: Data_out <= 16'h496C	;
				14'b00011000111010: Data_out <= 16'h4976	;
				14'b00011000111011: Data_out <= 16'h4980	;
				14'b00011000111100: Data_out <= 16'h498A	;
				14'b00011000111101: Data_out <= 16'h4995	;
				14'b00011000111110: Data_out <= 16'h499F	;
				14'b00011000111111: Data_out <= 16'h49A9	;
				14'b00011001000000: Data_out <= 16'h49B4	;
				14'b00011001000001: Data_out <= 16'h49BE	;
				14'b00011001000010: Data_out <= 16'h49C8	;
				14'b00011001000011: Data_out <= 16'h49D2	;
				14'b00011001000100: Data_out <= 16'h49DD	;
				14'b00011001000101: Data_out <= 16'h49E7	;
				14'b00011001000110: Data_out <= 16'h49F1	;
				14'b00011001000111: Data_out <= 16'h49FB	;
				14'b00011001001000: Data_out <= 16'h4A06	;
				14'b00011001001001: Data_out <= 16'h4A10	;
				14'b00011001001010: Data_out <= 16'h4A1A	;
				14'b00011001001011: Data_out <= 16'h4A24	;
				14'b00011001001100: Data_out <= 16'h4A2F	;
				14'b00011001001101: Data_out <= 16'h4A39	;
				14'b00011001001110: Data_out <= 16'h4A43	;
				14'b00011001001111: Data_out <= 16'h4A4D	;
				14'b00011001010000: Data_out <= 16'h4A58	;
				14'b00011001010001: Data_out <= 16'h4A62	;
				14'b00011001010010: Data_out <= 16'h4A6C	;
				14'b00011001010011: Data_out <= 16'h4A76	;
				14'b00011001010100: Data_out <= 16'h4A81	;
				14'b00011001010101: Data_out <= 16'h4A8B	;
				14'b00011001010110: Data_out <= 16'h4A95	;
				14'b00011001010111: Data_out <= 16'h4A9F	;
				14'b00011001011000: Data_out <= 16'h4AA9	;
				14'b00011001011001: Data_out <= 16'h4AB4	;
				14'b00011001011010: Data_out <= 16'h4ABE	;
				14'b00011001011011: Data_out <= 16'h4AC8	;
				14'b00011001011100: Data_out <= 16'h4AD2	;
				14'b00011001011101: Data_out <= 16'h4ADC	;
				14'b00011001011110: Data_out <= 16'h4AE7	;
				14'b00011001011111: Data_out <= 16'h4AF1	;
				14'b00011001100000: Data_out <= 16'h4AFB	;
				14'b00011001100001: Data_out <= 16'h4B05	;
				14'b00011001100010: Data_out <= 16'h4B0F	;
				14'b00011001100011: Data_out <= 16'h4B19	;
				14'b00011001100100: Data_out <= 16'h4B24	;
				14'b00011001100101: Data_out <= 16'h4B2E	;
				14'b00011001100110: Data_out <= 16'h4B38	;
				14'b00011001100111: Data_out <= 16'h4B42	;
				14'b00011001101000: Data_out <= 16'h4B4C	;
				14'b00011001101001: Data_out <= 16'h4B56	;
				14'b00011001101010: Data_out <= 16'h4B61	;
				14'b00011001101011: Data_out <= 16'h4B6B	;
				14'b00011001101100: Data_out <= 16'h4B75	;
				14'b00011001101101: Data_out <= 16'h4B7F	;
				14'b00011001101110: Data_out <= 16'h4B89	;
				14'b00011001101111: Data_out <= 16'h4B93	;
				14'b00011001110000: Data_out <= 16'h4B9E	;
				14'b00011001110001: Data_out <= 16'h4BA8	;
				14'b00011001110010: Data_out <= 16'h4BB2	;
				14'b00011001110011: Data_out <= 16'h4BBC	;
				14'b00011001110100: Data_out <= 16'h4BC6	;
				14'b00011001110101: Data_out <= 16'h4BD0	;
				14'b00011001110110: Data_out <= 16'h4BDA	;
				14'b00011001110111: Data_out <= 16'h4BE4	;
				14'b00011001111000: Data_out <= 16'h4BEF	;
				14'b00011001111001: Data_out <= 16'h4BF9	;
				14'b00011001111010: Data_out <= 16'h4C03	;
				14'b00011001111011: Data_out <= 16'h4C0D	;
				14'b00011001111100: Data_out <= 16'h4C17	;
				14'b00011001111101: Data_out <= 16'h4C21	;
				14'b00011001111110: Data_out <= 16'h4C2B	;
				14'b00011001111111: Data_out <= 16'h4C35	;
				14'b00011010000000: Data_out <= 16'h4C3F	;
				14'b00011010000001: Data_out <= 16'h4C49	;
				14'b00011010000010: Data_out <= 16'h4C54	;
				14'b00011010000011: Data_out <= 16'h4C5E	;
				14'b00011010000100: Data_out <= 16'h4C68	;
				14'b00011010000101: Data_out <= 16'h4C72	;
				14'b00011010000110: Data_out <= 16'h4C7C	;
				14'b00011010000111: Data_out <= 16'h4C86	;
				14'b00011010001000: Data_out <= 16'h4C90	;
				14'b00011010001001: Data_out <= 16'h4C9A	;
				14'b00011010001010: Data_out <= 16'h4CA4	;
				14'b00011010001011: Data_out <= 16'h4CAE	;
				14'b00011010001100: Data_out <= 16'h4CB8	;
				14'b00011010001101: Data_out <= 16'h4CC2	;
				14'b00011010001110: Data_out <= 16'h4CCC	;
				14'b00011010001111: Data_out <= 16'h4CD6	;
				14'b00011010010000: Data_out <= 16'h4CE1	;
				14'b00011010010001: Data_out <= 16'h4CEB	;
				14'b00011010010010: Data_out <= 16'h4CF5	;
				14'b00011010010011: Data_out <= 16'h4CFF	;
				14'b00011010010100: Data_out <= 16'h4D09	;
				14'b00011010010101: Data_out <= 16'h4D13	;
				14'b00011010010110: Data_out <= 16'h4D1D	;
				14'b00011010010111: Data_out <= 16'h4D27	;
				14'b00011010011000: Data_out <= 16'h4D31	;
				14'b00011010011001: Data_out <= 16'h4D3B	;
				14'b00011010011010: Data_out <= 16'h4D45	;
				14'b00011010011011: Data_out <= 16'h4D4F	;
				14'b00011010011100: Data_out <= 16'h4D59	;
				14'b00011010011101: Data_out <= 16'h4D63	;
				14'b00011010011110: Data_out <= 16'h4D6D	;
				14'b00011010011111: Data_out <= 16'h4D77	;
				14'b00011010100000: Data_out <= 16'h4D81	;
				14'b00011010100001: Data_out <= 16'h4D8B	;
				14'b00011010100010: Data_out <= 16'h4D95	;
				14'b00011010100011: Data_out <= 16'h4D9F	;
				14'b00011010100100: Data_out <= 16'h4DA9	;
				14'b00011010100101: Data_out <= 16'h4DB3	;
				14'b00011010100110: Data_out <= 16'h4DBD	;
				14'b00011010100111: Data_out <= 16'h4DC7	;
				14'b00011010101000: Data_out <= 16'h4DD1	;
				14'b00011010101001: Data_out <= 16'h4DDB	;
				14'b00011010101010: Data_out <= 16'h4DE5	;
				14'b00011010101011: Data_out <= 16'h4DEF	;
				14'b00011010101100: Data_out <= 16'h4DF9	;
				14'b00011010101101: Data_out <= 16'h4E03	;
				14'b00011010101110: Data_out <= 16'h4E0D	;
				14'b00011010101111: Data_out <= 16'h4E17	;
				14'b00011010110000: Data_out <= 16'h4E21	;
				14'b00011010110001: Data_out <= 16'h4E2A	;
				14'b00011010110010: Data_out <= 16'h4E34	;
				14'b00011010110011: Data_out <= 16'h4E3E	;
				14'b00011010110100: Data_out <= 16'h4E48	;
				14'b00011010110101: Data_out <= 16'h4E52	;
				14'b00011010110110: Data_out <= 16'h4E5C	;
				14'b00011010110111: Data_out <= 16'h4E66	;
				14'b00011010111000: Data_out <= 16'h4E70	;
				14'b00011010111001: Data_out <= 16'h4E7A	;
				14'b00011010111010: Data_out <= 16'h4E84	;
				14'b00011010111011: Data_out <= 16'h4E8E	;
				14'b00011010111100: Data_out <= 16'h4E98	;
				14'b00011010111101: Data_out <= 16'h4EA2	;
				14'b00011010111110: Data_out <= 16'h4EAC	;
				14'b00011010111111: Data_out <= 16'h4EB5	;
				14'b00011011000000: Data_out <= 16'h4EBF	;
				14'b00011011000001: Data_out <= 16'h4EC9	;
				14'b00011011000010: Data_out <= 16'h4ED3	;
				14'b00011011000011: Data_out <= 16'h4EDD	;
				14'b00011011000100: Data_out <= 16'h4EE7	;
				14'b00011011000101: Data_out <= 16'h4EF1	;
				14'b00011011000110: Data_out <= 16'h4EFB	;
				14'b00011011000111: Data_out <= 16'h4F05	;
				14'b00011011001000: Data_out <= 16'h4F0F	;
				14'b00011011001001: Data_out <= 16'h4F18	;
				14'b00011011001010: Data_out <= 16'h4F22	;
				14'b00011011001011: Data_out <= 16'h4F2C	;
				14'b00011011001100: Data_out <= 16'h4F36	;
				14'b00011011001101: Data_out <= 16'h4F40	;
				14'b00011011001110: Data_out <= 16'h4F4A	;
				14'b00011011001111: Data_out <= 16'h4F54	;
				14'b00011011010000: Data_out <= 16'h4F5E	;
				14'b00011011010001: Data_out <= 16'h4F67	;
				14'b00011011010010: Data_out <= 16'h4F71	;
				14'b00011011010011: Data_out <= 16'h4F7B	;
				14'b00011011010100: Data_out <= 16'h4F85	;
				14'b00011011010101: Data_out <= 16'h4F8F	;
				14'b00011011010110: Data_out <= 16'h4F99	;
				14'b00011011010111: Data_out <= 16'h4FA2	;
				14'b00011011011000: Data_out <= 16'h4FAC	;
				14'b00011011011001: Data_out <= 16'h4FB6	;
				14'b00011011011010: Data_out <= 16'h4FC0	;
				14'b00011011011011: Data_out <= 16'h4FCA	;
				14'b00011011011100: Data_out <= 16'h4FD4	;
				14'b00011011011101: Data_out <= 16'h4FDD	;
				14'b00011011011110: Data_out <= 16'h4FE7	;
				14'b00011011011111: Data_out <= 16'h4FF1	;
				14'b00011011100000: Data_out <= 16'h4FFB	;
				14'b00011011100001: Data_out <= 16'h5005	;
				14'b00011011100010: Data_out <= 16'h500E	;
				14'b00011011100011: Data_out <= 16'h5018	;
				14'b00011011100100: Data_out <= 16'h5022	;
				14'b00011011100101: Data_out <= 16'h502C	;
				14'b00011011100110: Data_out <= 16'h5036	;
				14'b00011011100111: Data_out <= 16'h503F	;
				14'b00011011101000: Data_out <= 16'h5049	;
				14'b00011011101001: Data_out <= 16'h5053	;
				14'b00011011101010: Data_out <= 16'h505D	;
				14'b00011011101011: Data_out <= 16'h5067	;
				14'b00011011101100: Data_out <= 16'h5070	;
				14'b00011011101101: Data_out <= 16'h507A	;
				14'b00011011101110: Data_out <= 16'h5084	;
				14'b00011011101111: Data_out <= 16'h508E	;
				14'b00011011110000: Data_out <= 16'h5097	;
				14'b00011011110001: Data_out <= 16'h50A1	;
				14'b00011011110010: Data_out <= 16'h50AB	;
				14'b00011011110011: Data_out <= 16'h50B5	;
				14'b00011011110100: Data_out <= 16'h50BE	;
				14'b00011011110101: Data_out <= 16'h50C8	;
				14'b00011011110110: Data_out <= 16'h50D2	;
				14'b00011011110111: Data_out <= 16'h50DC	;
				14'b00011011111000: Data_out <= 16'h50E5	;
				14'b00011011111001: Data_out <= 16'h50EF	;
				14'b00011011111010: Data_out <= 16'h50F9	;
				14'b00011011111011: Data_out <= 16'h5103	;
				14'b00011011111100: Data_out <= 16'h510C	;
				14'b00011011111101: Data_out <= 16'h5116	;
				14'b00011011111110: Data_out <= 16'h5120	;
				14'b00011011111111: Data_out <= 16'h512A	;
				14'b00011100000000: Data_out <= 16'h5133	;
				14'b00011100000001: Data_out <= 16'h513D	;
				14'b00011100000010: Data_out <= 16'h5147	;
				14'b00011100000011: Data_out <= 16'h5150	;
				14'b00011100000100: Data_out <= 16'h515A	;
				14'b00011100000101: Data_out <= 16'h5164	;
				14'b00011100000110: Data_out <= 16'h516D	;
				14'b00011100000111: Data_out <= 16'h5177	;
				14'b00011100001000: Data_out <= 16'h5181	;
				14'b00011100001001: Data_out <= 16'h518B	;
				14'b00011100001010: Data_out <= 16'h5194	;
				14'b00011100001011: Data_out <= 16'h519E	;
				14'b00011100001100: Data_out <= 16'h51A8	;
				14'b00011100001101: Data_out <= 16'h51B1	;
				14'b00011100001110: Data_out <= 16'h51BB	;
				14'b00011100001111: Data_out <= 16'h51C5	;
				14'b00011100010000: Data_out <= 16'h51CE	;
				14'b00011100010001: Data_out <= 16'h51D8	;
				14'b00011100010010: Data_out <= 16'h51E2	;
				14'b00011100010011: Data_out <= 16'h51EB	;
				14'b00011100010100: Data_out <= 16'h51F5	;
				14'b00011100010101: Data_out <= 16'h51FF	;
				14'b00011100010110: Data_out <= 16'h5208	;
				14'b00011100010111: Data_out <= 16'h5212	;
				14'b00011100011000: Data_out <= 16'h521C	;
				14'b00011100011001: Data_out <= 16'h5225	;
				14'b00011100011010: Data_out <= 16'h522F	;
				14'b00011100011011: Data_out <= 16'h5238	;
				14'b00011100011100: Data_out <= 16'h5242	;
				14'b00011100011101: Data_out <= 16'h524C	;
				14'b00011100011110: Data_out <= 16'h5255	;
				14'b00011100011111: Data_out <= 16'h525F	;
				14'b00011100100000: Data_out <= 16'h5269	;
				14'b00011100100001: Data_out <= 16'h5272	;
				14'b00011100100010: Data_out <= 16'h527C	;
				14'b00011100100011: Data_out <= 16'h5285	;
				14'b00011100100100: Data_out <= 16'h528F	;
				14'b00011100100101: Data_out <= 16'h5299	;
				14'b00011100100110: Data_out <= 16'h52A2	;
				14'b00011100100111: Data_out <= 16'h52AC	;
				14'b00011100101000: Data_out <= 16'h52B5	;
				14'b00011100101001: Data_out <= 16'h52BF	;
				14'b00011100101010: Data_out <= 16'h52C9	;
				14'b00011100101011: Data_out <= 16'h52D2	;
				14'b00011100101100: Data_out <= 16'h52DC	;
				14'b00011100101101: Data_out <= 16'h52E5	;
				14'b00011100101110: Data_out <= 16'h52EF	;
				14'b00011100101111: Data_out <= 16'h52F8	;
				14'b00011100110000: Data_out <= 16'h5302	;
				14'b00011100110001: Data_out <= 16'h530C	;
				14'b00011100110010: Data_out <= 16'h5315	;
				14'b00011100110011: Data_out <= 16'h531F	;
				14'b00011100110100: Data_out <= 16'h5328	;
				14'b00011100110101: Data_out <= 16'h5332	;
				14'b00011100110110: Data_out <= 16'h533B	;
				14'b00011100110111: Data_out <= 16'h5345	;
				14'b00011100111000: Data_out <= 16'h534E	;
				14'b00011100111001: Data_out <= 16'h5358	;
				14'b00011100111010: Data_out <= 16'h5361	;
				14'b00011100111011: Data_out <= 16'h536B	;
				14'b00011100111100: Data_out <= 16'h5375	;
				14'b00011100111101: Data_out <= 16'h537E	;
				14'b00011100111110: Data_out <= 16'h5388	;
				14'b00011100111111: Data_out <= 16'h5391	;
				14'b00011101000000: Data_out <= 16'h539B	;
				14'b00011101000001: Data_out <= 16'h53A4	;
				14'b00011101000010: Data_out <= 16'h53AE	;
				14'b00011101000011: Data_out <= 16'h53B7	;
				14'b00011101000100: Data_out <= 16'h53C1	;
				14'b00011101000101: Data_out <= 16'h53CA	;
				14'b00011101000110: Data_out <= 16'h53D4	;
				14'b00011101000111: Data_out <= 16'h53DD	;
				14'b00011101001000: Data_out <= 16'h53E7	;
				14'b00011101001001: Data_out <= 16'h53F0	;
				14'b00011101001010: Data_out <= 16'h53FA	;
				14'b00011101001011: Data_out <= 16'h5403	;
				14'b00011101001100: Data_out <= 16'h540D	;
				14'b00011101001101: Data_out <= 16'h5416	;
				14'b00011101001110: Data_out <= 16'h5420	;
				14'b00011101001111: Data_out <= 16'h5429	;
				14'b00011101010000: Data_out <= 16'h5432	;
				14'b00011101010001: Data_out <= 16'h543C	;
				14'b00011101010010: Data_out <= 16'h5445	;
				14'b00011101010011: Data_out <= 16'h544F	;
				14'b00011101010100: Data_out <= 16'h5458	;
				14'b00011101010101: Data_out <= 16'h5462	;
				14'b00011101010110: Data_out <= 16'h546B	;
				14'b00011101010111: Data_out <= 16'h5475	;
				14'b00011101011000: Data_out <= 16'h547E	;
				14'b00011101011001: Data_out <= 16'h5488	;
				14'b00011101011010: Data_out <= 16'h5491	;
				14'b00011101011011: Data_out <= 16'h549A	;
				14'b00011101011100: Data_out <= 16'h54A4	;
				14'b00011101011101: Data_out <= 16'h54AD	;
				14'b00011101011110: Data_out <= 16'h54B7	;
				14'b00011101011111: Data_out <= 16'h54C0	;
				14'b00011101100000: Data_out <= 16'h54C9	;
				14'b00011101100001: Data_out <= 16'h54D3	;
				14'b00011101100010: Data_out <= 16'h54DC	;
				14'b00011101100011: Data_out <= 16'h54E6	;
				14'b00011101100100: Data_out <= 16'h54EF	;
				14'b00011101100101: Data_out <= 16'h54F9	;
				14'b00011101100110: Data_out <= 16'h5502	;
				14'b00011101100111: Data_out <= 16'h550B	;
				14'b00011101101000: Data_out <= 16'h5515	;
				14'b00011101101001: Data_out <= 16'h551E	;
				14'b00011101101010: Data_out <= 16'h5527	;
				14'b00011101101011: Data_out <= 16'h5531	;
				14'b00011101101100: Data_out <= 16'h553A	;
				14'b00011101101101: Data_out <= 16'h5544	;
				14'b00011101101110: Data_out <= 16'h554D	;
				14'b00011101101111: Data_out <= 16'h5556	;
				14'b00011101110000: Data_out <= 16'h5560	;
				14'b00011101110001: Data_out <= 16'h5569	;
				14'b00011101110010: Data_out <= 16'h5572	;
				14'b00011101110011: Data_out <= 16'h557C	;
				14'b00011101110100: Data_out <= 16'h5585	;
				14'b00011101110101: Data_out <= 16'h558E	;
				14'b00011101110110: Data_out <= 16'h5598	;
				14'b00011101110111: Data_out <= 16'h55A1	;
				14'b00011101111000: Data_out <= 16'h55AA	;
				14'b00011101111001: Data_out <= 16'h55B4	;
				14'b00011101111010: Data_out <= 16'h55BD	;
				14'b00011101111011: Data_out <= 16'h55C6	;
				14'b00011101111100: Data_out <= 16'h55D0	;
				14'b00011101111101: Data_out <= 16'h55D9	;
				14'b00011101111110: Data_out <= 16'h55E2	;
				14'b00011101111111: Data_out <= 16'h55EC	;
				14'b00011110000000: Data_out <= 16'h55F5	;
				14'b00011110000001: Data_out <= 16'h55FE	;
				14'b00011110000010: Data_out <= 16'h5608	;
				14'b00011110000011: Data_out <= 16'h5611	;
				14'b00011110000100: Data_out <= 16'h561A	;
				14'b00011110000101: Data_out <= 16'h5624	;
				14'b00011110000110: Data_out <= 16'h562D	;
				14'b00011110000111: Data_out <= 16'h5636	;
				14'b00011110001000: Data_out <= 16'h563F	;
				14'b00011110001001: Data_out <= 16'h5649	;
				14'b00011110001010: Data_out <= 16'h5652	;
				14'b00011110001011: Data_out <= 16'h565B	;
				14'b00011110001100: Data_out <= 16'h5665	;
				14'b00011110001101: Data_out <= 16'h566E	;
				14'b00011110001110: Data_out <= 16'h5677	;
				14'b00011110001111: Data_out <= 16'h5680	;
				14'b00011110010000: Data_out <= 16'h568A	;
				14'b00011110010001: Data_out <= 16'h5693	;
				14'b00011110010010: Data_out <= 16'h569C	;
				14'b00011110010011: Data_out <= 16'h56A5	;
				14'b00011110010100: Data_out <= 16'h56AF	;
				14'b00011110010101: Data_out <= 16'h56B8	;
				14'b00011110010110: Data_out <= 16'h56C1	;
				14'b00011110010111: Data_out <= 16'h56CA	;
				14'b00011110011000: Data_out <= 16'h56D4	;
				14'b00011110011001: Data_out <= 16'h56DD	;
				14'b00011110011010: Data_out <= 16'h56E6	;
				14'b00011110011011: Data_out <= 16'h56EF	;
				14'b00011110011100: Data_out <= 16'h56F9	;
				14'b00011110011101: Data_out <= 16'h5702	;
				14'b00011110011110: Data_out <= 16'h570B	;
				14'b00011110011111: Data_out <= 16'h5714	;
				14'b00011110100000: Data_out <= 16'h571D	;
				14'b00011110100001: Data_out <= 16'h5727	;
				14'b00011110100010: Data_out <= 16'h5730	;
				14'b00011110100011: Data_out <= 16'h5739	;
				14'b00011110100100: Data_out <= 16'h5742	;
				14'b00011110100101: Data_out <= 16'h574B	;
				14'b00011110100110: Data_out <= 16'h5755	;
				14'b00011110100111: Data_out <= 16'h575E	;
				14'b00011110101000: Data_out <= 16'h5767	;
				14'b00011110101001: Data_out <= 16'h5770	;
				14'b00011110101010: Data_out <= 16'h5779	;
				14'b00011110101011: Data_out <= 16'h5782	;
				14'b00011110101100: Data_out <= 16'h578C	;
				14'b00011110101101: Data_out <= 16'h5795	;
				14'b00011110101110: Data_out <= 16'h579E	;
				14'b00011110101111: Data_out <= 16'h57A7	;
				14'b00011110110000: Data_out <= 16'h57B0	;
				14'b00011110110001: Data_out <= 16'h57B9	;
				14'b00011110110010: Data_out <= 16'h57C3	;
				14'b00011110110011: Data_out <= 16'h57CC	;
				14'b00011110110100: Data_out <= 16'h57D5	;
				14'b00011110110101: Data_out <= 16'h57DE	;
				14'b00011110110110: Data_out <= 16'h57E7	;
				14'b00011110110111: Data_out <= 16'h57F0	;
				14'b00011110111000: Data_out <= 16'h57F9	;
				14'b00011110111001: Data_out <= 16'h5802	;
				14'b00011110111010: Data_out <= 16'h580C	;
				14'b00011110111011: Data_out <= 16'h5815	;
				14'b00011110111100: Data_out <= 16'h581E	;
				14'b00011110111101: Data_out <= 16'h5827	;
				14'b00011110111110: Data_out <= 16'h5830	;
				14'b00011110111111: Data_out <= 16'h5839	;
				14'b00011111000000: Data_out <= 16'h5842	;
				14'b00011111000001: Data_out <= 16'h584B	;
				14'b00011111000010: Data_out <= 16'h5854	;
				14'b00011111000011: Data_out <= 16'h585E	;
				14'b00011111000100: Data_out <= 16'h5867	;
				14'b00011111000101: Data_out <= 16'h5870	;
				14'b00011111000110: Data_out <= 16'h5879	;
				14'b00011111000111: Data_out <= 16'h5882	;
				14'b00011111001000: Data_out <= 16'h588B	;
				14'b00011111001001: Data_out <= 16'h5894	;
				14'b00011111001010: Data_out <= 16'h589D	;
				14'b00011111001011: Data_out <= 16'h58A6	;
				14'b00011111001100: Data_out <= 16'h58AF	;
				14'b00011111001101: Data_out <= 16'h58B8	;
				14'b00011111001110: Data_out <= 16'h58C1	;
				14'b00011111001111: Data_out <= 16'h58CA	;
				14'b00011111010000: Data_out <= 16'h58D3	;
				14'b00011111010001: Data_out <= 16'h58DD	;
				14'b00011111010010: Data_out <= 16'h58E6	;
				14'b00011111010011: Data_out <= 16'h58EF	;
				14'b00011111010100: Data_out <= 16'h58F8	;
				14'b00011111010101: Data_out <= 16'h5901	;
				14'b00011111010110: Data_out <= 16'h590A	;
				14'b00011111010111: Data_out <= 16'h5913	;
				14'b00011111011000: Data_out <= 16'h591C	;
				14'b00011111011001: Data_out <= 16'h5925	;
				14'b00011111011010: Data_out <= 16'h592E	;
				14'b00011111011011: Data_out <= 16'h5937	;
				14'b00011111011100: Data_out <= 16'h5940	;
				14'b00011111011101: Data_out <= 16'h5949	;
				14'b00011111011110: Data_out <= 16'h5952	;
				14'b00011111011111: Data_out <= 16'h595B	;
				14'b00011111100000: Data_out <= 16'h5964	;
				14'b00011111100001: Data_out <= 16'h596D	;
				14'b00011111100010: Data_out <= 16'h5976	;
				14'b00011111100011: Data_out <= 16'h597F	;
				14'b00011111100100: Data_out <= 16'h5988	;
				14'b00011111100101: Data_out <= 16'h5991	;
				14'b00011111100110: Data_out <= 16'h599A	;
				14'b00011111100111: Data_out <= 16'h59A3	;
				14'b00011111101000: Data_out <= 16'h59AC	;
				14'b00011111101001: Data_out <= 16'h59B5	;
				14'b00011111101010: Data_out <= 16'h59BE	;
				14'b00011111101011: Data_out <= 16'h59C7	;
				14'b00011111101100: Data_out <= 16'h59CF	;
				14'b00011111101101: Data_out <= 16'h59D8	;
				14'b00011111101110: Data_out <= 16'h59E1	;
				14'b00011111101111: Data_out <= 16'h59EA	;
				14'b00011111110000: Data_out <= 16'h59F3	;
				14'b00011111110001: Data_out <= 16'h59FC	;
				14'b00011111110010: Data_out <= 16'h5A05	;
				14'b00011111110011: Data_out <= 16'h5A0E	;
				14'b00011111110100: Data_out <= 16'h5A17	;
				14'b00011111110101: Data_out <= 16'h5A20	;
				14'b00011111110110: Data_out <= 16'h5A29	;
				14'b00011111110111: Data_out <= 16'h5A32	;
				14'b00011111111000: Data_out <= 16'h5A3B	;
				14'b00011111111001: Data_out <= 16'h5A44	;
				14'b00011111111010: Data_out <= 16'h5A4C	;
				14'b00011111111011: Data_out <= 16'h5A55	;
				14'b00011111111100: Data_out <= 16'h5A5E	;
				14'b00011111111101: Data_out <= 16'h5A67	;
				14'b00011111111110: Data_out <= 16'h5A70	;
				14'b00011111111111: Data_out <= 16'h5A79	;
				14'b00100000000000: Data_out <= 16'h5A82	;
				14'b00100000000001: Data_out <= 16'h5A8B	;
				14'b00100000000010: Data_out <= 16'h5A94	;
				14'b00100000000011: Data_out <= 16'h5A9D	;
				14'b00100000000100: Data_out <= 16'h5AA5	;
				14'b00100000000101: Data_out <= 16'h5AAE	;
				14'b00100000000110: Data_out <= 16'h5AB7	;
				14'b00100000000111: Data_out <= 16'h5AC0	;
				14'b00100000001000: Data_out <= 16'h5AC9	;
				14'b00100000001001: Data_out <= 16'h5AD2	;
				14'b00100000001010: Data_out <= 16'h5ADB	;
				14'b00100000001011: Data_out <= 16'h5AE3	;
				14'b00100000001100: Data_out <= 16'h5AEC	;
				14'b00100000001101: Data_out <= 16'h5AF5	;
				14'b00100000001110: Data_out <= 16'h5AFE	;
				14'b00100000001111: Data_out <= 16'h5B07	;
				14'b00100000010000: Data_out <= 16'h5B10	;
				14'b00100000010001: Data_out <= 16'h5B18	;
				14'b00100000010010: Data_out <= 16'h5B21	;
				14'b00100000010011: Data_out <= 16'h5B2A	;
				14'b00100000010100: Data_out <= 16'h5B33	;
				14'b00100000010101: Data_out <= 16'h5B3C	;
				14'b00100000010110: Data_out <= 16'h5B45	;
				14'b00100000010111: Data_out <= 16'h5B4D	;
				14'b00100000011000: Data_out <= 16'h5B56	;
				14'b00100000011001: Data_out <= 16'h5B5F	;
				14'b00100000011010: Data_out <= 16'h5B68	;
				14'b00100000011011: Data_out <= 16'h5B71	;
				14'b00100000011100: Data_out <= 16'h5B79	;
				14'b00100000011101: Data_out <= 16'h5B82	;
				14'b00100000011110: Data_out <= 16'h5B8B	;
				14'b00100000011111: Data_out <= 16'h5B94	;
				14'b00100000100000: Data_out <= 16'h5B9C	;
				14'b00100000100001: Data_out <= 16'h5BA5	;
				14'b00100000100010: Data_out <= 16'h5BAE	;
				14'b00100000100011: Data_out <= 16'h5BB7	;
				14'b00100000100100: Data_out <= 16'h5BC0	;
				14'b00100000100101: Data_out <= 16'h5BC8	;
				14'b00100000100110: Data_out <= 16'h5BD1	;
				14'b00100000100111: Data_out <= 16'h5BDA	;
				14'b00100000101000: Data_out <= 16'h5BE3	;
				14'b00100000101001: Data_out <= 16'h5BEB	;
				14'b00100000101010: Data_out <= 16'h5BF4	;
				14'b00100000101011: Data_out <= 16'h5BFD	;
				14'b00100000101100: Data_out <= 16'h5C06	;
				14'b00100000101101: Data_out <= 16'h5C0E	;
				14'b00100000101110: Data_out <= 16'h5C17	;
				14'b00100000101111: Data_out <= 16'h5C20	;
				14'b00100000110000: Data_out <= 16'h5C28	;
				14'b00100000110001: Data_out <= 16'h5C31	;
				14'b00100000110010: Data_out <= 16'h5C3A	;
				14'b00100000110011: Data_out <= 16'h5C43	;
				14'b00100000110100: Data_out <= 16'h5C4B	;
				14'b00100000110101: Data_out <= 16'h5C54	;
				14'b00100000110110: Data_out <= 16'h5C5D	;
				14'b00100000110111: Data_out <= 16'h5C65	;
				14'b00100000111000: Data_out <= 16'h5C6E	;
				14'b00100000111001: Data_out <= 16'h5C77	;
				14'b00100000111010: Data_out <= 16'h5C7F	;
				14'b00100000111011: Data_out <= 16'h5C88	;
				14'b00100000111100: Data_out <= 16'h5C91	;
				14'b00100000111101: Data_out <= 16'h5C99	;
				14'b00100000111110: Data_out <= 16'h5CA2	;
				14'b00100000111111: Data_out <= 16'h5CAB	;
				14'b00100001000000: Data_out <= 16'h5CB4	;
				14'b00100001000001: Data_out <= 16'h5CBC	;
				14'b00100001000010: Data_out <= 16'h5CC5	;
				14'b00100001000011: Data_out <= 16'h5CCD	;
				14'b00100001000100: Data_out <= 16'h5CD6	;
				14'b00100001000101: Data_out <= 16'h5CDF	;
				14'b00100001000110: Data_out <= 16'h5CE7	;
				14'b00100001000111: Data_out <= 16'h5CF0	;
				14'b00100001001000: Data_out <= 16'h5CF9	;
				14'b00100001001001: Data_out <= 16'h5D01	;
				14'b00100001001010: Data_out <= 16'h5D0A	;
				14'b00100001001011: Data_out <= 16'h5D13	;
				14'b00100001001100: Data_out <= 16'h5D1B	;
				14'b00100001001101: Data_out <= 16'h5D24	;
				14'b00100001001110: Data_out <= 16'h5D2C	;
				14'b00100001001111: Data_out <= 16'h5D35	;
				14'b00100001010000: Data_out <= 16'h5D3E	;
				14'b00100001010001: Data_out <= 16'h5D46	;
				14'b00100001010010: Data_out <= 16'h5D4F	;
				14'b00100001010011: Data_out <= 16'h5D58	;
				14'b00100001010100: Data_out <= 16'h5D60	;
				14'b00100001010101: Data_out <= 16'h5D69	;
				14'b00100001010110: Data_out <= 16'h5D71	;
				14'b00100001010111: Data_out <= 16'h5D7A	;
				14'b00100001011000: Data_out <= 16'h5D82	;
				14'b00100001011001: Data_out <= 16'h5D8B	;
				14'b00100001011010: Data_out <= 16'h5D94	;
				14'b00100001011011: Data_out <= 16'h5D9C	;
				14'b00100001011100: Data_out <= 16'h5DA5	;
				14'b00100001011101: Data_out <= 16'h5DAD	;
				14'b00100001011110: Data_out <= 16'h5DB6	;
				14'b00100001011111: Data_out <= 16'h5DBE	;
				14'b00100001100000: Data_out <= 16'h5DC7	;
				14'b00100001100001: Data_out <= 16'h5DD0	;
				14'b00100001100010: Data_out <= 16'h5DD8	;
				14'b00100001100011: Data_out <= 16'h5DE1	;
				14'b00100001100100: Data_out <= 16'h5DE9	;
				14'b00100001100101: Data_out <= 16'h5DF2	;
				14'b00100001100110: Data_out <= 16'h5DFA	;
				14'b00100001100111: Data_out <= 16'h5E03	;
				14'b00100001101000: Data_out <= 16'h5E0B	;
				14'b00100001101001: Data_out <= 16'h5E14	;
				14'b00100001101010: Data_out <= 16'h5E1C	;
				14'b00100001101011: Data_out <= 16'h5E25	;
				14'b00100001101100: Data_out <= 16'h5E2D	;
				14'b00100001101101: Data_out <= 16'h5E36	;
				14'b00100001101110: Data_out <= 16'h5E3E	;
				14'b00100001101111: Data_out <= 16'h5E47	;
				14'b00100001110000: Data_out <= 16'h5E4F	;
				14'b00100001110001: Data_out <= 16'h5E58	;
				14'b00100001110010: Data_out <= 16'h5E60	;
				14'b00100001110011: Data_out <= 16'h5E69	;
				14'b00100001110100: Data_out <= 16'h5E71	;
				14'b00100001110101: Data_out <= 16'h5E7A	;
				14'b00100001110110: Data_out <= 16'h5E82	;
				14'b00100001110111: Data_out <= 16'h5E8B	;
				14'b00100001111000: Data_out <= 16'h5E93	;
				14'b00100001111001: Data_out <= 16'h5E9C	;
				14'b00100001111010: Data_out <= 16'h5EA4	;
				14'b00100001111011: Data_out <= 16'h5EAD	;
				14'b00100001111100: Data_out <= 16'h5EB5	;
				14'b00100001111101: Data_out <= 16'h5EBE	;
				14'b00100001111110: Data_out <= 16'h5EC6	;
				14'b00100001111111: Data_out <= 16'h5ECE	;
				14'b00100010000000: Data_out <= 16'h5ED7	;
				14'b00100010000001: Data_out <= 16'h5EDF	;
				14'b00100010000010: Data_out <= 16'h5EE8	;
				14'b00100010000011: Data_out <= 16'h5EF0	;
				14'b00100010000100: Data_out <= 16'h5EF9	;
				14'b00100010000101: Data_out <= 16'h5F01	;
				14'b00100010000110: Data_out <= 16'h5F09	;
				14'b00100010000111: Data_out <= 16'h5F12	;
				14'b00100010001000: Data_out <= 16'h5F1A	;
				14'b00100010001001: Data_out <= 16'h5F23	;
				14'b00100010001010: Data_out <= 16'h5F2B	;
				14'b00100010001011: Data_out <= 16'h5F33	;
				14'b00100010001100: Data_out <= 16'h5F3C	;
				14'b00100010001101: Data_out <= 16'h5F44	;
				14'b00100010001110: Data_out <= 16'h5F4D	;
				14'b00100010001111: Data_out <= 16'h5F55	;
				14'b00100010010000: Data_out <= 16'h5F5D	;
				14'b00100010010001: Data_out <= 16'h5F66	;
				14'b00100010010010: Data_out <= 16'h5F6E	;
				14'b00100010010011: Data_out <= 16'h5F77	;
				14'b00100010010100: Data_out <= 16'h5F7F	;
				14'b00100010010101: Data_out <= 16'h5F87	;
				14'b00100010010110: Data_out <= 16'h5F90	;
				14'b00100010010111: Data_out <= 16'h5F98	;
				14'b00100010011000: Data_out <= 16'h5FA0	;
				14'b00100010011001: Data_out <= 16'h5FA9	;
				14'b00100010011010: Data_out <= 16'h5FB1	;
				14'b00100010011011: Data_out <= 16'h5FB9	;
				14'b00100010011100: Data_out <= 16'h5FC2	;
				14'b00100010011101: Data_out <= 16'h5FCA	;
				14'b00100010011110: Data_out <= 16'h5FD2	;
				14'b00100010011111: Data_out <= 16'h5FDB	;
				14'b00100010100000: Data_out <= 16'h5FE3	;
				14'b00100010100001: Data_out <= 16'h5FEB	;
				14'b00100010100010: Data_out <= 16'h5FF4	;
				14'b00100010100011: Data_out <= 16'h5FFC	;
				14'b00100010100100: Data_out <= 16'h6004	;
				14'b00100010100101: Data_out <= 16'h600D	;
				14'b00100010100110: Data_out <= 16'h6015	;
				14'b00100010100111: Data_out <= 16'h601D	;
				14'b00100010101000: Data_out <= 16'h6026	;
				14'b00100010101001: Data_out <= 16'h602E	;
				14'b00100010101010: Data_out <= 16'h6036	;
				14'b00100010101011: Data_out <= 16'h603E	;
				14'b00100010101100: Data_out <= 16'h6047	;
				14'b00100010101101: Data_out <= 16'h604F	;
				14'b00100010101110: Data_out <= 16'h6057	;
				14'b00100010101111: Data_out <= 16'h6060	;
				14'b00100010110000: Data_out <= 16'h6068	;
				14'b00100010110001: Data_out <= 16'h6070	;
				14'b00100010110010: Data_out <= 16'h6078	;
				14'b00100010110011: Data_out <= 16'h6081	;
				14'b00100010110100: Data_out <= 16'h6089	;
				14'b00100010110101: Data_out <= 16'h6091	;
				14'b00100010110110: Data_out <= 16'h6099	;
				14'b00100010110111: Data_out <= 16'h60A2	;
				14'b00100010111000: Data_out <= 16'h60AA	;
				14'b00100010111001: Data_out <= 16'h60B2	;
				14'b00100010111010: Data_out <= 16'h60BA	;
				14'b00100010111011: Data_out <= 16'h60C2	;
				14'b00100010111100: Data_out <= 16'h60CB	;
				14'b00100010111101: Data_out <= 16'h60D3	;
				14'b00100010111110: Data_out <= 16'h60DB	;
				14'b00100010111111: Data_out <= 16'h60E3	;
				14'b00100011000000: Data_out <= 16'h60EC	;
				14'b00100011000001: Data_out <= 16'h60F4	;
				14'b00100011000010: Data_out <= 16'h60FC	;
				14'b00100011000011: Data_out <= 16'h6104	;
				14'b00100011000100: Data_out <= 16'h610C	;
				14'b00100011000101: Data_out <= 16'h6115	;
				14'b00100011000110: Data_out <= 16'h611D	;
				14'b00100011000111: Data_out <= 16'h6125	;
				14'b00100011001000: Data_out <= 16'h612D	;
				14'b00100011001001: Data_out <= 16'h6135	;
				14'b00100011001010: Data_out <= 16'h613D	;
				14'b00100011001011: Data_out <= 16'h6146	;
				14'b00100011001100: Data_out <= 16'h614E	;
				14'b00100011001101: Data_out <= 16'h6156	;
				14'b00100011001110: Data_out <= 16'h615E	;
				14'b00100011001111: Data_out <= 16'h6166	;
				14'b00100011010000: Data_out <= 16'h616E	;
				14'b00100011010001: Data_out <= 16'h6177	;
				14'b00100011010010: Data_out <= 16'h617F	;
				14'b00100011010011: Data_out <= 16'h6187	;
				14'b00100011010100: Data_out <= 16'h618F	;
				14'b00100011010101: Data_out <= 16'h6197	;
				14'b00100011010110: Data_out <= 16'h619F	;
				14'b00100011010111: Data_out <= 16'h61A7	;
				14'b00100011011000: Data_out <= 16'h61AF	;
				14'b00100011011001: Data_out <= 16'h61B8	;
				14'b00100011011010: Data_out <= 16'h61C0	;
				14'b00100011011011: Data_out <= 16'h61C8	;
				14'b00100011011100: Data_out <= 16'h61D0	;
				14'b00100011011101: Data_out <= 16'h61D8	;
				14'b00100011011110: Data_out <= 16'h61E0	;
				14'b00100011011111: Data_out <= 16'h61E8	;
				14'b00100011100000: Data_out <= 16'h61F0	;
				14'b00100011100001: Data_out <= 16'h61F8	;
				14'b00100011100010: Data_out <= 16'h6201	;
				14'b00100011100011: Data_out <= 16'h6209	;
				14'b00100011100100: Data_out <= 16'h6211	;
				14'b00100011100101: Data_out <= 16'h6219	;
				14'b00100011100110: Data_out <= 16'h6221	;
				14'b00100011100111: Data_out <= 16'h6229	;
				14'b00100011101000: Data_out <= 16'h6231	;
				14'b00100011101001: Data_out <= 16'h6239	;
				14'b00100011101010: Data_out <= 16'h6241	;
				14'b00100011101011: Data_out <= 16'h6249	;
				14'b00100011101100: Data_out <= 16'h6251	;
				14'b00100011101101: Data_out <= 16'h6259	;
				14'b00100011101110: Data_out <= 16'h6261	;
				14'b00100011101111: Data_out <= 16'h6269	;
				14'b00100011110000: Data_out <= 16'h6271	;
				14'b00100011110001: Data_out <= 16'h6279	;
				14'b00100011110010: Data_out <= 16'h6281	;
				14'b00100011110011: Data_out <= 16'h6289	;
				14'b00100011110100: Data_out <= 16'h6291	;
				14'b00100011110101: Data_out <= 16'h6299	;
				14'b00100011110110: Data_out <= 16'h62A1	;
				14'b00100011110111: Data_out <= 16'h62A9	;
				14'b00100011111000: Data_out <= 16'h62B1	;
				14'b00100011111001: Data_out <= 16'h62B9	;
				14'b00100011111010: Data_out <= 16'h62C1	;
				14'b00100011111011: Data_out <= 16'h62C9	;
				14'b00100011111100: Data_out <= 16'h62D1	;
				14'b00100011111101: Data_out <= 16'h62D9	;
				14'b00100011111110: Data_out <= 16'h62E1	;
				14'b00100011111111: Data_out <= 16'h62E9	;
				14'b00100100000000: Data_out <= 16'h62F1	;
				14'b00100100000001: Data_out <= 16'h62F9	;
				14'b00100100000010: Data_out <= 16'h6301	;
				14'b00100100000011: Data_out <= 16'h6309	;
				14'b00100100000100: Data_out <= 16'h6311	;
				14'b00100100000101: Data_out <= 16'h6319	;
				14'b00100100000110: Data_out <= 16'h6321	;
				14'b00100100000111: Data_out <= 16'h6329	;
				14'b00100100001000: Data_out <= 16'h6331	;
				14'b00100100001001: Data_out <= 16'h6339	;
				14'b00100100001010: Data_out <= 16'h6341	;
				14'b00100100001011: Data_out <= 16'h6349	;
				14'b00100100001100: Data_out <= 16'h6351	;
				14'b00100100001101: Data_out <= 16'h6359	;
				14'b00100100001110: Data_out <= 16'h6361	;
				14'b00100100001111: Data_out <= 16'h6368	;
				14'b00100100010000: Data_out <= 16'h6370	;
				14'b00100100010001: Data_out <= 16'h6378	;
				14'b00100100010010: Data_out <= 16'h6380	;
				14'b00100100010011: Data_out <= 16'h6388	;
				14'b00100100010100: Data_out <= 16'h6390	;
				14'b00100100010101: Data_out <= 16'h6398	;
				14'b00100100010110: Data_out <= 16'h63A0	;
				14'b00100100010111: Data_out <= 16'h63A8	;
				14'b00100100011000: Data_out <= 16'h63B0	;
				14'b00100100011001: Data_out <= 16'h63B7	;
				14'b00100100011010: Data_out <= 16'h63BF	;
				14'b00100100011011: Data_out <= 16'h63C7	;
				14'b00100100011100: Data_out <= 16'h63CF	;
				14'b00100100011101: Data_out <= 16'h63D7	;
				14'b00100100011110: Data_out <= 16'h63DF	;
				14'b00100100011111: Data_out <= 16'h63E7	;
				14'b00100100100000: Data_out <= 16'h63EF	;
				14'b00100100100001: Data_out <= 16'h63F6	;
				14'b00100100100010: Data_out <= 16'h63FE	;
				14'b00100100100011: Data_out <= 16'h6406	;
				14'b00100100100100: Data_out <= 16'h640E	;
				14'b00100100100101: Data_out <= 16'h6416	;
				14'b00100100100110: Data_out <= 16'h641E	;
				14'b00100100100111: Data_out <= 16'h6425	;
				14'b00100100101000: Data_out <= 16'h642D	;
				14'b00100100101001: Data_out <= 16'h6435	;
				14'b00100100101010: Data_out <= 16'h643D	;
				14'b00100100101011: Data_out <= 16'h6445	;
				14'b00100100101100: Data_out <= 16'h644C	;
				14'b00100100101101: Data_out <= 16'h6454	;
				14'b00100100101110: Data_out <= 16'h645C	;
				14'b00100100101111: Data_out <= 16'h6464	;
				14'b00100100110000: Data_out <= 16'h646C	;
				14'b00100100110001: Data_out <= 16'h6473	;
				14'b00100100110010: Data_out <= 16'h647B	;
				14'b00100100110011: Data_out <= 16'h6483	;
				14'b00100100110100: Data_out <= 16'h648B	;
				14'b00100100110101: Data_out <= 16'h6493	;
				14'b00100100110110: Data_out <= 16'h649A	;
				14'b00100100110111: Data_out <= 16'h64A2	;
				14'b00100100111000: Data_out <= 16'h64AA	;
				14'b00100100111001: Data_out <= 16'h64B2	;
				14'b00100100111010: Data_out <= 16'h64B9	;
				14'b00100100111011: Data_out <= 16'h64C1	;
				14'b00100100111100: Data_out <= 16'h64C9	;
				14'b00100100111101: Data_out <= 16'h64D1	;
				14'b00100100111110: Data_out <= 16'h64D8	;
				14'b00100100111111: Data_out <= 16'h64E0	;
				14'b00100101000000: Data_out <= 16'h64E8	;
				14'b00100101000001: Data_out <= 16'h64F0	;
				14'b00100101000010: Data_out <= 16'h64F7	;
				14'b00100101000011: Data_out <= 16'h64FF	;
				14'b00100101000100: Data_out <= 16'h6507	;
				14'b00100101000101: Data_out <= 16'h650E	;
				14'b00100101000110: Data_out <= 16'h6516	;
				14'b00100101000111: Data_out <= 16'h651E	;
				14'b00100101001000: Data_out <= 16'h6526	;
				14'b00100101001001: Data_out <= 16'h652D	;
				14'b00100101001010: Data_out <= 16'h6535	;
				14'b00100101001011: Data_out <= 16'h653D	;
				14'b00100101001100: Data_out <= 16'h6544	;
				14'b00100101001101: Data_out <= 16'h654C	;
				14'b00100101001110: Data_out <= 16'h6554	;
				14'b00100101001111: Data_out <= 16'h655B	;
				14'b00100101010000: Data_out <= 16'h6563	;
				14'b00100101010001: Data_out <= 16'h656B	;
				14'b00100101010010: Data_out <= 16'h6572	;
				14'b00100101010011: Data_out <= 16'h657A	;
				14'b00100101010100: Data_out <= 16'h6582	;
				14'b00100101010101: Data_out <= 16'h6589	;
				14'b00100101010110: Data_out <= 16'h6591	;
				14'b00100101010111: Data_out <= 16'h6599	;
				14'b00100101011000: Data_out <= 16'h65A0	;
				14'b00100101011001: Data_out <= 16'h65A8	;
				14'b00100101011010: Data_out <= 16'h65B0	;
				14'b00100101011011: Data_out <= 16'h65B7	;
				14'b00100101011100: Data_out <= 16'h65BF	;
				14'b00100101011101: Data_out <= 16'h65C6	;
				14'b00100101011110: Data_out <= 16'h65CE	;
				14'b00100101011111: Data_out <= 16'h65D6	;
				14'b00100101100000: Data_out <= 16'h65DD	;
				14'b00100101100001: Data_out <= 16'h65E5	;
				14'b00100101100010: Data_out <= 16'h65EC	;
				14'b00100101100011: Data_out <= 16'h65F4	;
				14'b00100101100100: Data_out <= 16'h65FC	;
				14'b00100101100101: Data_out <= 16'h6603	;
				14'b00100101100110: Data_out <= 16'h660B	;
				14'b00100101100111: Data_out <= 16'h6612	;
				14'b00100101101000: Data_out <= 16'h661A	;
				14'b00100101101001: Data_out <= 16'h6622	;
				14'b00100101101010: Data_out <= 16'h6629	;
				14'b00100101101011: Data_out <= 16'h6631	;
				14'b00100101101100: Data_out <= 16'h6638	;
				14'b00100101101101: Data_out <= 16'h6640	;
				14'b00100101101110: Data_out <= 16'h6647	;
				14'b00100101101111: Data_out <= 16'h664F	;
				14'b00100101110000: Data_out <= 16'h6657	;
				14'b00100101110001: Data_out <= 16'h665E	;
				14'b00100101110010: Data_out <= 16'h6666	;
				14'b00100101110011: Data_out <= 16'h666D	;
				14'b00100101110100: Data_out <= 16'h6675	;
				14'b00100101110101: Data_out <= 16'h667C	;
				14'b00100101110110: Data_out <= 16'h6684	;
				14'b00100101110111: Data_out <= 16'h668B	;
				14'b00100101111000: Data_out <= 16'h6693	;
				14'b00100101111001: Data_out <= 16'h669A	;
				14'b00100101111010: Data_out <= 16'h66A2	;
				14'b00100101111011: Data_out <= 16'h66A9	;
				14'b00100101111100: Data_out <= 16'h66B1	;
				14'b00100101111101: Data_out <= 16'h66B8	;
				14'b00100101111110: Data_out <= 16'h66C0	;
				14'b00100101111111: Data_out <= 16'h66C7	;
				14'b00100110000000: Data_out <= 16'h66CF	;
				14'b00100110000001: Data_out <= 16'h66D6	;
				14'b00100110000010: Data_out <= 16'h66DE	;
				14'b00100110000011: Data_out <= 16'h66E5	;
				14'b00100110000100: Data_out <= 16'h66ED	;
				14'b00100110000101: Data_out <= 16'h66F4	;
				14'b00100110000110: Data_out <= 16'h66FC	;
				14'b00100110000111: Data_out <= 16'h6703	;
				14'b00100110001000: Data_out <= 16'h670B	;
				14'b00100110001001: Data_out <= 16'h6712	;
				14'b00100110001010: Data_out <= 16'h6719	;
				14'b00100110001011: Data_out <= 16'h6721	;
				14'b00100110001100: Data_out <= 16'h6728	;
				14'b00100110001101: Data_out <= 16'h6730	;
				14'b00100110001110: Data_out <= 16'h6737	;
				14'b00100110001111: Data_out <= 16'h673F	;
				14'b00100110010000: Data_out <= 16'h6746	;
				14'b00100110010001: Data_out <= 16'h674D	;
				14'b00100110010010: Data_out <= 16'h6755	;
				14'b00100110010011: Data_out <= 16'h675C	;
				14'b00100110010100: Data_out <= 16'h6764	;
				14'b00100110010101: Data_out <= 16'h676B	;
				14'b00100110010110: Data_out <= 16'h6773	;
				14'b00100110010111: Data_out <= 16'h677A	;
				14'b00100110011000: Data_out <= 16'h6781	;
				14'b00100110011001: Data_out <= 16'h6789	;
				14'b00100110011010: Data_out <= 16'h6790	;
				14'b00100110011011: Data_out <= 16'h6797	;
				14'b00100110011100: Data_out <= 16'h679F	;
				14'b00100110011101: Data_out <= 16'h67A6	;
				14'b00100110011110: Data_out <= 16'h67AE	;
				14'b00100110011111: Data_out <= 16'h67B5	;
				14'b00100110100000: Data_out <= 16'h67BC	;
				14'b00100110100001: Data_out <= 16'h67C4	;
				14'b00100110100010: Data_out <= 16'h67CB	;
				14'b00100110100011: Data_out <= 16'h67D2	;
				14'b00100110100100: Data_out <= 16'h67DA	;
				14'b00100110100101: Data_out <= 16'h67E1	;
				14'b00100110100110: Data_out <= 16'h67E8	;
				14'b00100110100111: Data_out <= 16'h67F0	;
				14'b00100110101000: Data_out <= 16'h67F7	;
				14'b00100110101001: Data_out <= 16'h67FE	;
				14'b00100110101010: Data_out <= 16'h6806	;
				14'b00100110101011: Data_out <= 16'h680D	;
				14'b00100110101100: Data_out <= 16'h6814	;
				14'b00100110101101: Data_out <= 16'h681C	;
				14'b00100110101110: Data_out <= 16'h6823	;
				14'b00100110101111: Data_out <= 16'h682A	;
				14'b00100110110000: Data_out <= 16'h6832	;
				14'b00100110110001: Data_out <= 16'h6839	;
				14'b00100110110010: Data_out <= 16'h6840	;
				14'b00100110110011: Data_out <= 16'h6848	;
				14'b00100110110100: Data_out <= 16'h684F	;
				14'b00100110110101: Data_out <= 16'h6856	;
				14'b00100110110110: Data_out <= 16'h685D	;
				14'b00100110110111: Data_out <= 16'h6865	;
				14'b00100110111000: Data_out <= 16'h686C	;
				14'b00100110111001: Data_out <= 16'h6873	;
				14'b00100110111010: Data_out <= 16'h687A	;
				14'b00100110111011: Data_out <= 16'h6882	;
				14'b00100110111100: Data_out <= 16'h6889	;
				14'b00100110111101: Data_out <= 16'h6890	;
				14'b00100110111110: Data_out <= 16'h6897	;
				14'b00100110111111: Data_out <= 16'h689F	;
				14'b00100111000000: Data_out <= 16'h68A6	;
				14'b00100111000001: Data_out <= 16'h68AD	;
				14'b00100111000010: Data_out <= 16'h68B4	;
				14'b00100111000011: Data_out <= 16'h68BC	;
				14'b00100111000100: Data_out <= 16'h68C3	;
				14'b00100111000101: Data_out <= 16'h68CA	;
				14'b00100111000110: Data_out <= 16'h68D1	;
				14'b00100111000111: Data_out <= 16'h68D8	;
				14'b00100111001000: Data_out <= 16'h68E0	;
				14'b00100111001001: Data_out <= 16'h68E7	;
				14'b00100111001010: Data_out <= 16'h68EE	;
				14'b00100111001011: Data_out <= 16'h68F5	;
				14'b00100111001100: Data_out <= 16'h68FC	;
				14'b00100111001101: Data_out <= 16'h6904	;
				14'b00100111001110: Data_out <= 16'h690B	;
				14'b00100111001111: Data_out <= 16'h6912	;
				14'b00100111010000: Data_out <= 16'h6919	;
				14'b00100111010001: Data_out <= 16'h6920	;
				14'b00100111010010: Data_out <= 16'h6928	;
				14'b00100111010011: Data_out <= 16'h692F	;
				14'b00100111010100: Data_out <= 16'h6936	;
				14'b00100111010101: Data_out <= 16'h693D	;
				14'b00100111010110: Data_out <= 16'h6944	;
				14'b00100111010111: Data_out <= 16'h694B	;
				14'b00100111011000: Data_out <= 16'h6952	;
				14'b00100111011001: Data_out <= 16'h695A	;
				14'b00100111011010: Data_out <= 16'h6961	;
				14'b00100111011011: Data_out <= 16'h6968	;
				14'b00100111011100: Data_out <= 16'h696F	;
				14'b00100111011101: Data_out <= 16'h6976	;
				14'b00100111011110: Data_out <= 16'h697D	;
				14'b00100111011111: Data_out <= 16'h6984	;
				14'b00100111100000: Data_out <= 16'h698B	;
				14'b00100111100001: Data_out <= 16'h6993	;
				14'b00100111100010: Data_out <= 16'h699A	;
				14'b00100111100011: Data_out <= 16'h69A1	;
				14'b00100111100100: Data_out <= 16'h69A8	;
				14'b00100111100101: Data_out <= 16'h69AF	;
				14'b00100111100110: Data_out <= 16'h69B6	;
				14'b00100111100111: Data_out <= 16'h69BD	;
				14'b00100111101000: Data_out <= 16'h69C4	;
				14'b00100111101001: Data_out <= 16'h69CB	;
				14'b00100111101010: Data_out <= 16'h69D2	;
				14'b00100111101011: Data_out <= 16'h69D9	;
				14'b00100111101100: Data_out <= 16'h69E0	;
				14'b00100111101101: Data_out <= 16'h69E7	;
				14'b00100111101110: Data_out <= 16'h69EF	;
				14'b00100111101111: Data_out <= 16'h69F6	;
				14'b00100111110000: Data_out <= 16'h69FD	;
				14'b00100111110001: Data_out <= 16'h6A04	;
				14'b00100111110010: Data_out <= 16'h6A0B	;
				14'b00100111110011: Data_out <= 16'h6A12	;
				14'b00100111110100: Data_out <= 16'h6A19	;
				14'b00100111110101: Data_out <= 16'h6A20	;
				14'b00100111110110: Data_out <= 16'h6A27	;
				14'b00100111110111: Data_out <= 16'h6A2E	;
				14'b00100111111000: Data_out <= 16'h6A35	;
				14'b00100111111001: Data_out <= 16'h6A3C	;
				14'b00100111111010: Data_out <= 16'h6A43	;
				14'b00100111111011: Data_out <= 16'h6A4A	;
				14'b00100111111100: Data_out <= 16'h6A51	;
				14'b00100111111101: Data_out <= 16'h6A58	;
				14'b00100111111110: Data_out <= 16'h6A5F	;
				14'b00100111111111: Data_out <= 16'h6A66	;
				14'b00101000000000: Data_out <= 16'h6A6D	;
				14'b00101000000001: Data_out <= 16'h6A74	;
				14'b00101000000010: Data_out <= 16'h6A7B	;
				14'b00101000000011: Data_out <= 16'h6A82	;
				14'b00101000000100: Data_out <= 16'h6A89	;
				14'b00101000000101: Data_out <= 16'h6A90	;
				14'b00101000000110: Data_out <= 16'h6A97	;
				14'b00101000000111: Data_out <= 16'h6A9E	;
				14'b00101000001000: Data_out <= 16'h6AA5	;
				14'b00101000001001: Data_out <= 16'h6AAC	;
				14'b00101000001010: Data_out <= 16'h6AB2	;
				14'b00101000001011: Data_out <= 16'h6AB9	;
				14'b00101000001100: Data_out <= 16'h6AC0	;
				14'b00101000001101: Data_out <= 16'h6AC7	;
				14'b00101000001110: Data_out <= 16'h6ACE	;
				14'b00101000001111: Data_out <= 16'h6AD5	;
				14'b00101000010000: Data_out <= 16'h6ADC	;
				14'b00101000010001: Data_out <= 16'h6AE3	;
				14'b00101000010010: Data_out <= 16'h6AEA	;
				14'b00101000010011: Data_out <= 16'h6AF1	;
				14'b00101000010100: Data_out <= 16'h6AF8	;
				14'b00101000010101: Data_out <= 16'h6AFF	;
				14'b00101000010110: Data_out <= 16'h6B05	;
				14'b00101000010111: Data_out <= 16'h6B0C	;
				14'b00101000011000: Data_out <= 16'h6B13	;
				14'b00101000011001: Data_out <= 16'h6B1A	;
				14'b00101000011010: Data_out <= 16'h6B21	;
				14'b00101000011011: Data_out <= 16'h6B28	;
				14'b00101000011100: Data_out <= 16'h6B2F	;
				14'b00101000011101: Data_out <= 16'h6B36	;
				14'b00101000011110: Data_out <= 16'h6B3C	;
				14'b00101000011111: Data_out <= 16'h6B43	;
				14'b00101000100000: Data_out <= 16'h6B4A	;
				14'b00101000100001: Data_out <= 16'h6B51	;
				14'b00101000100010: Data_out <= 16'h6B58	;
				14'b00101000100011: Data_out <= 16'h6B5F	;
				14'b00101000100100: Data_out <= 16'h6B66	;
				14'b00101000100101: Data_out <= 16'h6B6C	;
				14'b00101000100110: Data_out <= 16'h6B73	;
				14'b00101000100111: Data_out <= 16'h6B7A	;
				14'b00101000101000: Data_out <= 16'h6B81	;
				14'b00101000101001: Data_out <= 16'h6B88	;
				14'b00101000101010: Data_out <= 16'h6B8F	;
				14'b00101000101011: Data_out <= 16'h6B95	;
				14'b00101000101100: Data_out <= 16'h6B9C	;
				14'b00101000101101: Data_out <= 16'h6BA3	;
				14'b00101000101110: Data_out <= 16'h6BAA	;
				14'b00101000101111: Data_out <= 16'h6BB1	;
				14'b00101000110000: Data_out <= 16'h6BB7	;
				14'b00101000110001: Data_out <= 16'h6BBE	;
				14'b00101000110010: Data_out <= 16'h6BC5	;
				14'b00101000110011: Data_out <= 16'h6BCC	;
				14'b00101000110100: Data_out <= 16'h6BD2	;
				14'b00101000110101: Data_out <= 16'h6BD9	;
				14'b00101000110110: Data_out <= 16'h6BE0	;
				14'b00101000110111: Data_out <= 16'h6BE7	;
				14'b00101000111000: Data_out <= 16'h6BEE	;
				14'b00101000111001: Data_out <= 16'h6BF4	;
				14'b00101000111010: Data_out <= 16'h6BFB	;
				14'b00101000111011: Data_out <= 16'h6C02	;
				14'b00101000111100: Data_out <= 16'h6C08	;
				14'b00101000111101: Data_out <= 16'h6C0F	;
				14'b00101000111110: Data_out <= 16'h6C16	;
				14'b00101000111111: Data_out <= 16'h6C1D	;
				14'b00101001000000: Data_out <= 16'h6C23	;
				14'b00101001000001: Data_out <= 16'h6C2A	;
				14'b00101001000010: Data_out <= 16'h6C31	;
				14'b00101001000011: Data_out <= 16'h6C38	;
				14'b00101001000100: Data_out <= 16'h6C3E	;
				14'b00101001000101: Data_out <= 16'h6C45	;
				14'b00101001000110: Data_out <= 16'h6C4C	;
				14'b00101001000111: Data_out <= 16'h6C52	;
				14'b00101001001000: Data_out <= 16'h6C59	;
				14'b00101001001001: Data_out <= 16'h6C60	;
				14'b00101001001010: Data_out <= 16'h6C66	;
				14'b00101001001011: Data_out <= 16'h6C6D	;
				14'b00101001001100: Data_out <= 16'h6C74	;
				14'b00101001001101: Data_out <= 16'h6C7A	;
				14'b00101001001110: Data_out <= 16'h6C81	;
				14'b00101001001111: Data_out <= 16'h6C88	;
				14'b00101001010000: Data_out <= 16'h6C8E	;
				14'b00101001010001: Data_out <= 16'h6C95	;
				14'b00101001010010: Data_out <= 16'h6C9C	;
				14'b00101001010011: Data_out <= 16'h6CA2	;
				14'b00101001010100: Data_out <= 16'h6CA9	;
				14'b00101001010101: Data_out <= 16'h6CB0	;
				14'b00101001010110: Data_out <= 16'h6CB6	;
				14'b00101001010111: Data_out <= 16'h6CBD	;
				14'b00101001011000: Data_out <= 16'h6CC4	;
				14'b00101001011001: Data_out <= 16'h6CCA	;
				14'b00101001011010: Data_out <= 16'h6CD1	;
				14'b00101001011011: Data_out <= 16'h6CD7	;
				14'b00101001011100: Data_out <= 16'h6CDE	;
				14'b00101001011101: Data_out <= 16'h6CE5	;
				14'b00101001011110: Data_out <= 16'h6CEB	;
				14'b00101001011111: Data_out <= 16'h6CF2	;
				14'b00101001100000: Data_out <= 16'h6CF8	;
				14'b00101001100001: Data_out <= 16'h6CFF	;
				14'b00101001100010: Data_out <= 16'h6D06	;
				14'b00101001100011: Data_out <= 16'h6D0C	;
				14'b00101001100100: Data_out <= 16'h6D13	;
				14'b00101001100101: Data_out <= 16'h6D19	;
				14'b00101001100110: Data_out <= 16'h6D20	;
				14'b00101001100111: Data_out <= 16'h6D26	;
				14'b00101001101000: Data_out <= 16'h6D2D	;
				14'b00101001101001: Data_out <= 16'h6D34	;
				14'b00101001101010: Data_out <= 16'h6D3A	;
				14'b00101001101011: Data_out <= 16'h6D41	;
				14'b00101001101100: Data_out <= 16'h6D47	;
				14'b00101001101101: Data_out <= 16'h6D4E	;
				14'b00101001101110: Data_out <= 16'h6D54	;
				14'b00101001101111: Data_out <= 16'h6D5B	;
				14'b00101001110000: Data_out <= 16'h6D61	;
				14'b00101001110001: Data_out <= 16'h6D68	;
				14'b00101001110010: Data_out <= 16'h6D6E	;
				14'b00101001110011: Data_out <= 16'h6D75	;
				14'b00101001110100: Data_out <= 16'h6D7B	;
				14'b00101001110101: Data_out <= 16'h6D82	;
				14'b00101001110110: Data_out <= 16'h6D88	;
				14'b00101001110111: Data_out <= 16'h6D8F	;
				14'b00101001111000: Data_out <= 16'h6D95	;
				14'b00101001111001: Data_out <= 16'h6D9C	;
				14'b00101001111010: Data_out <= 16'h6DA2	;
				14'b00101001111011: Data_out <= 16'h6DA9	;
				14'b00101001111100: Data_out <= 16'h6DAF	;
				14'b00101001111101: Data_out <= 16'h6DB6	;
				14'b00101001111110: Data_out <= 16'h6DBC	;
				14'b00101001111111: Data_out <= 16'h6DC3	;
				14'b00101010000000: Data_out <= 16'h6DC9	;
				14'b00101010000001: Data_out <= 16'h6DD0	;
				14'b00101010000010: Data_out <= 16'h6DD6	;
				14'b00101010000011: Data_out <= 16'h6DDD	;
				14'b00101010000100: Data_out <= 16'h6DE3	;
				14'b00101010000101: Data_out <= 16'h6DEA	;
				14'b00101010000110: Data_out <= 16'h6DF0	;
				14'b00101010000111: Data_out <= 16'h6DF6	;
				14'b00101010001000: Data_out <= 16'h6DFD	;
				14'b00101010001001: Data_out <= 16'h6E03	;
				14'b00101010001010: Data_out <= 16'h6E0A	;
				14'b00101010001011: Data_out <= 16'h6E10	;
				14'b00101010001100: Data_out <= 16'h6E17	;
				14'b00101010001101: Data_out <= 16'h6E1D	;
				14'b00101010001110: Data_out <= 16'h6E23	;
				14'b00101010001111: Data_out <= 16'h6E2A	;
				14'b00101010010000: Data_out <= 16'h6E30	;
				14'b00101010010001: Data_out <= 16'h6E37	;
				14'b00101010010010: Data_out <= 16'h6E3D	;
				14'b00101010010011: Data_out <= 16'h6E43	;
				14'b00101010010100: Data_out <= 16'h6E4A	;
				14'b00101010010101: Data_out <= 16'h6E50	;
				14'b00101010010110: Data_out <= 16'h6E56	;
				14'b00101010010111: Data_out <= 16'h6E5D	;
				14'b00101010011000: Data_out <= 16'h6E63	;
				14'b00101010011001: Data_out <= 16'h6E6A	;
				14'b00101010011010: Data_out <= 16'h6E70	;
				14'b00101010011011: Data_out <= 16'h6E76	;
				14'b00101010011100: Data_out <= 16'h6E7D	;
				14'b00101010011101: Data_out <= 16'h6E83	;
				14'b00101010011110: Data_out <= 16'h6E89	;
				14'b00101010011111: Data_out <= 16'h6E90	;
				14'b00101010100000: Data_out <= 16'h6E96	;
				14'b00101010100001: Data_out <= 16'h6E9C	;
				14'b00101010100010: Data_out <= 16'h6EA3	;
				14'b00101010100011: Data_out <= 16'h6EA9	;
				14'b00101010100100: Data_out <= 16'h6EAF	;
				14'b00101010100101: Data_out <= 16'h6EB5	;
				14'b00101010100110: Data_out <= 16'h6EBC	;
				14'b00101010100111: Data_out <= 16'h6EC2	;
				14'b00101010101000: Data_out <= 16'h6EC8	;
				14'b00101010101001: Data_out <= 16'h6ECF	;
				14'b00101010101010: Data_out <= 16'h6ED5	;
				14'b00101010101011: Data_out <= 16'h6EDB	;
				14'b00101010101100: Data_out <= 16'h6EE2	;
				14'b00101010101101: Data_out <= 16'h6EE8	;
				14'b00101010101110: Data_out <= 16'h6EEE	;
				14'b00101010101111: Data_out <= 16'h6EF4	;
				14'b00101010110000: Data_out <= 16'h6EFB	;
				14'b00101010110001: Data_out <= 16'h6F01	;
				14'b00101010110010: Data_out <= 16'h6F07	;
				14'b00101010110011: Data_out <= 16'h6F0D	;
				14'b00101010110100: Data_out <= 16'h6F14	;
				14'b00101010110101: Data_out <= 16'h6F1A	;
				14'b00101010110110: Data_out <= 16'h6F20	;
				14'b00101010110111: Data_out <= 16'h6F26	;
				14'b00101010111000: Data_out <= 16'h6F2D	;
				14'b00101010111001: Data_out <= 16'h6F33	;
				14'b00101010111010: Data_out <= 16'h6F39	;
				14'b00101010111011: Data_out <= 16'h6F3F	;
				14'b00101010111100: Data_out <= 16'h6F45	;
				14'b00101010111101: Data_out <= 16'h6F4C	;
				14'b00101010111110: Data_out <= 16'h6F52	;
				14'b00101010111111: Data_out <= 16'h6F58	;
				14'b00101011000000: Data_out <= 16'h6F5E	;
				14'b00101011000001: Data_out <= 16'h6F64	;
				14'b00101011000010: Data_out <= 16'h6F6B	;
				14'b00101011000011: Data_out <= 16'h6F71	;
				14'b00101011000100: Data_out <= 16'h6F77	;
				14'b00101011000101: Data_out <= 16'h6F7D	;
				14'b00101011000110: Data_out <= 16'h6F83	;
				14'b00101011000111: Data_out <= 16'h6F89	;
				14'b00101011001000: Data_out <= 16'h6F90	;
				14'b00101011001001: Data_out <= 16'h6F96	;
				14'b00101011001010: Data_out <= 16'h6F9C	;
				14'b00101011001011: Data_out <= 16'h6FA2	;
				14'b00101011001100: Data_out <= 16'h6FA8	;
				14'b00101011001101: Data_out <= 16'h6FAE	;
				14'b00101011001110: Data_out <= 16'h6FB5	;
				14'b00101011001111: Data_out <= 16'h6FBB	;
				14'b00101011010000: Data_out <= 16'h6FC1	;
				14'b00101011010001: Data_out <= 16'h6FC7	;
				14'b00101011010010: Data_out <= 16'h6FCD	;
				14'b00101011010011: Data_out <= 16'h6FD3	;
				14'b00101011010100: Data_out <= 16'h6FD9	;
				14'b00101011010101: Data_out <= 16'h6FDF	;
				14'b00101011010110: Data_out <= 16'h6FE5	;
				14'b00101011010111: Data_out <= 16'h6FEC	;
				14'b00101011011000: Data_out <= 16'h6FF2	;
				14'b00101011011001: Data_out <= 16'h6FF8	;
				14'b00101011011010: Data_out <= 16'h6FFE	;
				14'b00101011011011: Data_out <= 16'h7004	;
				14'b00101011011100: Data_out <= 16'h700A	;
				14'b00101011011101: Data_out <= 16'h7010	;
				14'b00101011011110: Data_out <= 16'h7016	;
				14'b00101011011111: Data_out <= 16'h701C	;
				14'b00101011100000: Data_out <= 16'h7022	;
				14'b00101011100001: Data_out <= 16'h7028	;
				14'b00101011100010: Data_out <= 16'h702E	;
				14'b00101011100011: Data_out <= 16'h7034	;
				14'b00101011100100: Data_out <= 16'h703A	;
				14'b00101011100101: Data_out <= 16'h7041	;
				14'b00101011100110: Data_out <= 16'h7047	;
				14'b00101011100111: Data_out <= 16'h704D	;
				14'b00101011101000: Data_out <= 16'h7053	;
				14'b00101011101001: Data_out <= 16'h7059	;
				14'b00101011101010: Data_out <= 16'h705F	;
				14'b00101011101011: Data_out <= 16'h7065	;
				14'b00101011101100: Data_out <= 16'h706B	;
				14'b00101011101101: Data_out <= 16'h7071	;
				14'b00101011101110: Data_out <= 16'h7077	;
				14'b00101011101111: Data_out <= 16'h707D	;
				14'b00101011110000: Data_out <= 16'h7083	;
				14'b00101011110001: Data_out <= 16'h7089	;
				14'b00101011110010: Data_out <= 16'h708F	;
				14'b00101011110011: Data_out <= 16'h7095	;
				14'b00101011110100: Data_out <= 16'h709B	;
				14'b00101011110101: Data_out <= 16'h70A1	;
				14'b00101011110110: Data_out <= 16'h70A7	;
				14'b00101011110111: Data_out <= 16'h70AD	;
				14'b00101011111000: Data_out <= 16'h70B2	;
				14'b00101011111001: Data_out <= 16'h70B8	;
				14'b00101011111010: Data_out <= 16'h70BE	;
				14'b00101011111011: Data_out <= 16'h70C4	;
				14'b00101011111100: Data_out <= 16'h70CA	;
				14'b00101011111101: Data_out <= 16'h70D0	;
				14'b00101011111110: Data_out <= 16'h70D6	;
				14'b00101011111111: Data_out <= 16'h70DC	;
				14'b00101100000000: Data_out <= 16'h70E2	;
				14'b00101100000001: Data_out <= 16'h70E8	;
				14'b00101100000010: Data_out <= 16'h70EE	;
				14'b00101100000011: Data_out <= 16'h70F4	;
				14'b00101100000100: Data_out <= 16'h70FA	;
				14'b00101100000101: Data_out <= 16'h7100	;
				14'b00101100000110: Data_out <= 16'h7105	;
				14'b00101100000111: Data_out <= 16'h710B	;
				14'b00101100001000: Data_out <= 16'h7111	;
				14'b00101100001001: Data_out <= 16'h7117	;
				14'b00101100001010: Data_out <= 16'h711D	;
				14'b00101100001011: Data_out <= 16'h7123	;
				14'b00101100001100: Data_out <= 16'h7129	;
				14'b00101100001101: Data_out <= 16'h712F	;
				14'b00101100001110: Data_out <= 16'h7135	;
				14'b00101100001111: Data_out <= 16'h713A	;
				14'b00101100010000: Data_out <= 16'h7140	;
				14'b00101100010001: Data_out <= 16'h7146	;
				14'b00101100010010: Data_out <= 16'h714C	;
				14'b00101100010011: Data_out <= 16'h7152	;
				14'b00101100010100: Data_out <= 16'h7158	;
				14'b00101100010101: Data_out <= 16'h715D	;
				14'b00101100010110: Data_out <= 16'h7163	;
				14'b00101100010111: Data_out <= 16'h7169	;
				14'b00101100011000: Data_out <= 16'h716F	;
				14'b00101100011001: Data_out <= 16'h7175	;
				14'b00101100011010: Data_out <= 16'h717B	;
				14'b00101100011011: Data_out <= 16'h7180	;
				14'b00101100011100: Data_out <= 16'h7186	;
				14'b00101100011101: Data_out <= 16'h718C	;
				14'b00101100011110: Data_out <= 16'h7192	;
				14'b00101100011111: Data_out <= 16'h7198	;
				14'b00101100100000: Data_out <= 16'h719D	;
				14'b00101100100001: Data_out <= 16'h71A3	;
				14'b00101100100010: Data_out <= 16'h71A9	;
				14'b00101100100011: Data_out <= 16'h71AF	;
				14'b00101100100100: Data_out <= 16'h71B5	;
				14'b00101100100101: Data_out <= 16'h71BA	;
				14'b00101100100110: Data_out <= 16'h71C0	;
				14'b00101100100111: Data_out <= 16'h71C6	;
				14'b00101100101000: Data_out <= 16'h71CC	;
				14'b00101100101001: Data_out <= 16'h71D1	;
				14'b00101100101010: Data_out <= 16'h71D7	;
				14'b00101100101011: Data_out <= 16'h71DD	;
				14'b00101100101100: Data_out <= 16'h71E3	;
				14'b00101100101101: Data_out <= 16'h71E8	;
				14'b00101100101110: Data_out <= 16'h71EE	;
				14'b00101100101111: Data_out <= 16'h71F4	;
				14'b00101100110000: Data_out <= 16'h71F9	;
				14'b00101100110001: Data_out <= 16'h71FF	;
				14'b00101100110010: Data_out <= 16'h7205	;
				14'b00101100110011: Data_out <= 16'h720B	;
				14'b00101100110100: Data_out <= 16'h7210	;
				14'b00101100110101: Data_out <= 16'h7216	;
				14'b00101100110110: Data_out <= 16'h721C	;
				14'b00101100110111: Data_out <= 16'h7221	;
				14'b00101100111000: Data_out <= 16'h7227	;
				14'b00101100111001: Data_out <= 16'h722D	;
				14'b00101100111010: Data_out <= 16'h7232	;
				14'b00101100111011: Data_out <= 16'h7238	;
				14'b00101100111100: Data_out <= 16'h723E	;
				14'b00101100111101: Data_out <= 16'h7243	;
				14'b00101100111110: Data_out <= 16'h7249	;
				14'b00101100111111: Data_out <= 16'h724F	;
				14'b00101101000000: Data_out <= 16'h7254	;
				14'b00101101000001: Data_out <= 16'h725A	;
				14'b00101101000010: Data_out <= 16'h7260	;
				14'b00101101000011: Data_out <= 16'h7265	;
				14'b00101101000100: Data_out <= 16'h726B	;
				14'b00101101000101: Data_out <= 16'h7271	;
				14'b00101101000110: Data_out <= 16'h7276	;
				14'b00101101000111: Data_out <= 16'h727C	;
				14'b00101101001000: Data_out <= 16'h7281	;
				14'b00101101001001: Data_out <= 16'h7287	;
				14'b00101101001010: Data_out <= 16'h728D	;
				14'b00101101001011: Data_out <= 16'h7292	;
				14'b00101101001100: Data_out <= 16'h7298	;
				14'b00101101001101: Data_out <= 16'h729D	;
				14'b00101101001110: Data_out <= 16'h72A3	;
				14'b00101101001111: Data_out <= 16'h72A9	;
				14'b00101101010000: Data_out <= 16'h72AE	;
				14'b00101101010001: Data_out <= 16'h72B4	;
				14'b00101101010010: Data_out <= 16'h72B9	;
				14'b00101101010011: Data_out <= 16'h72BF	;
				14'b00101101010100: Data_out <= 16'h72C5	;
				14'b00101101010101: Data_out <= 16'h72CA	;
				14'b00101101010110: Data_out <= 16'h72D0	;
				14'b00101101010111: Data_out <= 16'h72D5	;
				14'b00101101011000: Data_out <= 16'h72DB	;
				14'b00101101011001: Data_out <= 16'h72E0	;
				14'b00101101011010: Data_out <= 16'h72E6	;
				14'b00101101011011: Data_out <= 16'h72EB	;
				14'b00101101011100: Data_out <= 16'h72F1	;
				14'b00101101011101: Data_out <= 16'h72F6	;
				14'b00101101011110: Data_out <= 16'h72FC	;
				14'b00101101011111: Data_out <= 16'h7301	;
				14'b00101101100000: Data_out <= 16'h7307	;
				14'b00101101100001: Data_out <= 16'h730C	;
				14'b00101101100010: Data_out <= 16'h7312	;
				14'b00101101100011: Data_out <= 16'h7317	;
				14'b00101101100100: Data_out <= 16'h731D	;
				14'b00101101100101: Data_out <= 16'h7322	;
				14'b00101101100110: Data_out <= 16'h7328	;
				14'b00101101100111: Data_out <= 16'h732D	;
				14'b00101101101000: Data_out <= 16'h7333	;
				14'b00101101101001: Data_out <= 16'h7338	;
				14'b00101101101010: Data_out <= 16'h733E	;
				14'b00101101101011: Data_out <= 16'h7343	;
				14'b00101101101100: Data_out <= 16'h7349	;
				14'b00101101101101: Data_out <= 16'h734E	;
				14'b00101101101110: Data_out <= 16'h7354	;
				14'b00101101101111: Data_out <= 16'h7359	;
				14'b00101101110000: Data_out <= 16'h735F	;
				14'b00101101110001: Data_out <= 16'h7364	;
				14'b00101101110010: Data_out <= 16'h7369	;
				14'b00101101110011: Data_out <= 16'h736F	;
				14'b00101101110100: Data_out <= 16'h7374	;
				14'b00101101110101: Data_out <= 16'h737A	;
				14'b00101101110110: Data_out <= 16'h737F	;
				14'b00101101110111: Data_out <= 16'h7385	;
				14'b00101101111000: Data_out <= 16'h738A	;
				14'b00101101111001: Data_out <= 16'h738F	;
				14'b00101101111010: Data_out <= 16'h7395	;
				14'b00101101111011: Data_out <= 16'h739A	;
				14'b00101101111100: Data_out <= 16'h73A0	;
				14'b00101101111101: Data_out <= 16'h73A5	;
				14'b00101101111110: Data_out <= 16'h73AA	;
				14'b00101101111111: Data_out <= 16'h73B0	;
				14'b00101110000000: Data_out <= 16'h73B5	;
				14'b00101110000001: Data_out <= 16'h73BA	;
				14'b00101110000010: Data_out <= 16'h73C0	;
				14'b00101110000011: Data_out <= 16'h73C5	;
				14'b00101110000100: Data_out <= 16'h73CB	;
				14'b00101110000101: Data_out <= 16'h73D0	;
				14'b00101110000110: Data_out <= 16'h73D5	;
				14'b00101110000111: Data_out <= 16'h73DB	;
				14'b00101110001000: Data_out <= 16'h73E0	;
				14'b00101110001001: Data_out <= 16'h73E5	;
				14'b00101110001010: Data_out <= 16'h73EB	;
				14'b00101110001011: Data_out <= 16'h73F0	;
				14'b00101110001100: Data_out <= 16'h73F5	;
				14'b00101110001101: Data_out <= 16'h73FB	;
				14'b00101110001110: Data_out <= 16'h7400	;
				14'b00101110001111: Data_out <= 16'h7405	;
				14'b00101110010000: Data_out <= 16'h740B	;
				14'b00101110010001: Data_out <= 16'h7410	;
				14'b00101110010010: Data_out <= 16'h7415	;
				14'b00101110010011: Data_out <= 16'h741A	;
				14'b00101110010100: Data_out <= 16'h7420	;
				14'b00101110010101: Data_out <= 16'h7425	;
				14'b00101110010110: Data_out <= 16'h742A	;
				14'b00101110010111: Data_out <= 16'h7430	;
				14'b00101110011000: Data_out <= 16'h7435	;
				14'b00101110011001: Data_out <= 16'h743A	;
				14'b00101110011010: Data_out <= 16'h743F	;
				14'b00101110011011: Data_out <= 16'h7445	;
				14'b00101110011100: Data_out <= 16'h744A	;
				14'b00101110011101: Data_out <= 16'h744F	;
				14'b00101110011110: Data_out <= 16'h7454	;
				14'b00101110011111: Data_out <= 16'h745A	;
				14'b00101110100000: Data_out <= 16'h745F	;
				14'b00101110100001: Data_out <= 16'h7464	;
				14'b00101110100010: Data_out <= 16'h7469	;
				14'b00101110100011: Data_out <= 16'h746E	;
				14'b00101110100100: Data_out <= 16'h7474	;
				14'b00101110100101: Data_out <= 16'h7479	;
				14'b00101110100110: Data_out <= 16'h747E	;
				14'b00101110100111: Data_out <= 16'h7483	;
				14'b00101110101000: Data_out <= 16'h7489	;
				14'b00101110101001: Data_out <= 16'h748E	;
				14'b00101110101010: Data_out <= 16'h7493	;
				14'b00101110101011: Data_out <= 16'h7498	;
				14'b00101110101100: Data_out <= 16'h749D	;
				14'b00101110101101: Data_out <= 16'h74A2	;
				14'b00101110101110: Data_out <= 16'h74A8	;
				14'b00101110101111: Data_out <= 16'h74AD	;
				14'b00101110110000: Data_out <= 16'h74B2	;
				14'b00101110110001: Data_out <= 16'h74B7	;
				14'b00101110110010: Data_out <= 16'h74BC	;
				14'b00101110110011: Data_out <= 16'h74C1	;
				14'b00101110110100: Data_out <= 16'h74C7	;
				14'b00101110110101: Data_out <= 16'h74CC	;
				14'b00101110110110: Data_out <= 16'h74D1	;
				14'b00101110110111: Data_out <= 16'h74D6	;
				14'b00101110111000: Data_out <= 16'h74DB	;
				14'b00101110111001: Data_out <= 16'h74E0	;
				14'b00101110111010: Data_out <= 16'h74E5	;
				14'b00101110111011: Data_out <= 16'h74EA	;
				14'b00101110111100: Data_out <= 16'h74F0	;
				14'b00101110111101: Data_out <= 16'h74F5	;
				14'b00101110111110: Data_out <= 16'h74FA	;
				14'b00101110111111: Data_out <= 16'h74FF	;
				14'b00101111000000: Data_out <= 16'h7504	;
				14'b00101111000001: Data_out <= 16'h7509	;
				14'b00101111000010: Data_out <= 16'h750E	;
				14'b00101111000011: Data_out <= 16'h7513	;
				14'b00101111000100: Data_out <= 16'h7518	;
				14'b00101111000101: Data_out <= 16'h751D	;
				14'b00101111000110: Data_out <= 16'h7522	;
				14'b00101111000111: Data_out <= 16'h7528	;
				14'b00101111001000: Data_out <= 16'h752D	;
				14'b00101111001001: Data_out <= 16'h7532	;
				14'b00101111001010: Data_out <= 16'h7537	;
				14'b00101111001011: Data_out <= 16'h753C	;
				14'b00101111001100: Data_out <= 16'h7541	;
				14'b00101111001101: Data_out <= 16'h7546	;
				14'b00101111001110: Data_out <= 16'h754B	;
				14'b00101111001111: Data_out <= 16'h7550	;
				14'b00101111010000: Data_out <= 16'h7555	;
				14'b00101111010001: Data_out <= 16'h755A	;
				14'b00101111010010: Data_out <= 16'h755F	;
				14'b00101111010011: Data_out <= 16'h7564	;
				14'b00101111010100: Data_out <= 16'h7569	;
				14'b00101111010101: Data_out <= 16'h756E	;
				14'b00101111010110: Data_out <= 16'h7573	;
				14'b00101111010111: Data_out <= 16'h7578	;
				14'b00101111011000: Data_out <= 16'h757D	;
				14'b00101111011001: Data_out <= 16'h7582	;
				14'b00101111011010: Data_out <= 16'h7587	;
				14'b00101111011011: Data_out <= 16'h758C	;
				14'b00101111011100: Data_out <= 16'h7591	;
				14'b00101111011101: Data_out <= 16'h7596	;
				14'b00101111011110: Data_out <= 16'h759B	;
				14'b00101111011111: Data_out <= 16'h75A0	;
				14'b00101111100000: Data_out <= 16'h75A5	;
				14'b00101111100001: Data_out <= 16'h75AA	;
				14'b00101111100010: Data_out <= 16'h75AF	;
				14'b00101111100011: Data_out <= 16'h75B4	;
				14'b00101111100100: Data_out <= 16'h75B8	;
				14'b00101111100101: Data_out <= 16'h75BD	;
				14'b00101111100110: Data_out <= 16'h75C2	;
				14'b00101111100111: Data_out <= 16'h75C7	;
				14'b00101111101000: Data_out <= 16'h75CC	;
				14'b00101111101001: Data_out <= 16'h75D1	;
				14'b00101111101010: Data_out <= 16'h75D6	;
				14'b00101111101011: Data_out <= 16'h75DB	;
				14'b00101111101100: Data_out <= 16'h75E0	;
				14'b00101111101101: Data_out <= 16'h75E5	;
				14'b00101111101110: Data_out <= 16'h75EA	;
				14'b00101111101111: Data_out <= 16'h75EE	;
				14'b00101111110000: Data_out <= 16'h75F3	;
				14'b00101111110001: Data_out <= 16'h75F8	;
				14'b00101111110010: Data_out <= 16'h75FD	;
				14'b00101111110011: Data_out <= 16'h7602	;
				14'b00101111110100: Data_out <= 16'h7607	;
				14'b00101111110101: Data_out <= 16'h760C	;
				14'b00101111110110: Data_out <= 16'h7611	;
				14'b00101111110111: Data_out <= 16'h7615	;
				14'b00101111111000: Data_out <= 16'h761A	;
				14'b00101111111001: Data_out <= 16'h761F	;
				14'b00101111111010: Data_out <= 16'h7624	;
				14'b00101111111011: Data_out <= 16'h7629	;
				14'b00101111111100: Data_out <= 16'h762E	;
				14'b00101111111101: Data_out <= 16'h7632	;
				14'b00101111111110: Data_out <= 16'h7637	;
				14'b00101111111111: Data_out <= 16'h763C	;
				14'b00110000000000: Data_out <= 16'h7641	;
				14'b00110000000001: Data_out <= 16'h7646	;
				14'b00110000000010: Data_out <= 16'h764A	;
				14'b00110000000011: Data_out <= 16'h764F	;
				14'b00110000000100: Data_out <= 16'h7654	;
				14'b00110000000101: Data_out <= 16'h7659	;
				14'b00110000000110: Data_out <= 16'h765E	;
				14'b00110000000111: Data_out <= 16'h7662	;
				14'b00110000001000: Data_out <= 16'h7667	;
				14'b00110000001001: Data_out <= 16'h766C	;
				14'b00110000001010: Data_out <= 16'h7671	;
				14'b00110000001011: Data_out <= 16'h7675	;
				14'b00110000001100: Data_out <= 16'h767A	;
				14'b00110000001101: Data_out <= 16'h767F	;
				14'b00110000001110: Data_out <= 16'h7684	;
				14'b00110000001111: Data_out <= 16'h7688	;
				14'b00110000010000: Data_out <= 16'h768D	;
				14'b00110000010001: Data_out <= 16'h7692	;
				14'b00110000010010: Data_out <= 16'h7697	;
				14'b00110000010011: Data_out <= 16'h769B	;
				14'b00110000010100: Data_out <= 16'h76A0	;
				14'b00110000010101: Data_out <= 16'h76A5	;
				14'b00110000010110: Data_out <= 16'h76AA	;
				14'b00110000010111: Data_out <= 16'h76AE	;
				14'b00110000011000: Data_out <= 16'h76B3	;
				14'b00110000011001: Data_out <= 16'h76B8	;
				14'b00110000011010: Data_out <= 16'h76BC	;
				14'b00110000011011: Data_out <= 16'h76C1	;
				14'b00110000011100: Data_out <= 16'h76C6	;
				14'b00110000011101: Data_out <= 16'h76CA	;
				14'b00110000011110: Data_out <= 16'h76CF	;
				14'b00110000011111: Data_out <= 16'h76D4	;
				14'b00110000100000: Data_out <= 16'h76D8	;
				14'b00110000100001: Data_out <= 16'h76DD	;
				14'b00110000100010: Data_out <= 16'h76E2	;
				14'b00110000100011: Data_out <= 16'h76E6	;
				14'b00110000100100: Data_out <= 16'h76EB	;
				14'b00110000100101: Data_out <= 16'h76F0	;
				14'b00110000100110: Data_out <= 16'h76F4	;
				14'b00110000100111: Data_out <= 16'h76F9	;
				14'b00110000101000: Data_out <= 16'h76FE	;
				14'b00110000101001: Data_out <= 16'h7702	;
				14'b00110000101010: Data_out <= 16'h7707	;
				14'b00110000101011: Data_out <= 16'h770C	;
				14'b00110000101100: Data_out <= 16'h7710	;
				14'b00110000101101: Data_out <= 16'h7715	;
				14'b00110000101110: Data_out <= 16'h7719	;
				14'b00110000101111: Data_out <= 16'h771E	;
				14'b00110000110000: Data_out <= 16'h7723	;
				14'b00110000110001: Data_out <= 16'h7727	;
				14'b00110000110010: Data_out <= 16'h772C	;
				14'b00110000110011: Data_out <= 16'h7730	;
				14'b00110000110100: Data_out <= 16'h7735	;
				14'b00110000110101: Data_out <= 16'h7739	;
				14'b00110000110110: Data_out <= 16'h773E	;
				14'b00110000110111: Data_out <= 16'h7743	;
				14'b00110000111000: Data_out <= 16'h7747	;
				14'b00110000111001: Data_out <= 16'h774C	;
				14'b00110000111010: Data_out <= 16'h7750	;
				14'b00110000111011: Data_out <= 16'h7755	;
				14'b00110000111100: Data_out <= 16'h7759	;
				14'b00110000111101: Data_out <= 16'h775E	;
				14'b00110000111110: Data_out <= 16'h7762	;
				14'b00110000111111: Data_out <= 16'h7767	;
				14'b00110001000000: Data_out <= 16'h776B	;
				14'b00110001000001: Data_out <= 16'h7770	;
				14'b00110001000010: Data_out <= 16'h7775	;
				14'b00110001000011: Data_out <= 16'h7779	;
				14'b00110001000100: Data_out <= 16'h777E	;
				14'b00110001000101: Data_out <= 16'h7782	;
				14'b00110001000110: Data_out <= 16'h7787	;
				14'b00110001000111: Data_out <= 16'h778B	;
				14'b00110001001000: Data_out <= 16'h7790	;
				14'b00110001001001: Data_out <= 16'h7794	;
				14'b00110001001010: Data_out <= 16'h7798	;
				14'b00110001001011: Data_out <= 16'h779D	;
				14'b00110001001100: Data_out <= 16'h77A1	;
				14'b00110001001101: Data_out <= 16'h77A6	;
				14'b00110001001110: Data_out <= 16'h77AA	;
				14'b00110001001111: Data_out <= 16'h77AF	;
				14'b00110001010000: Data_out <= 16'h77B3	;
				14'b00110001010001: Data_out <= 16'h77B8	;
				14'b00110001010010: Data_out <= 16'h77BC	;
				14'b00110001010011: Data_out <= 16'h77C1	;
				14'b00110001010100: Data_out <= 16'h77C5	;
				14'b00110001010101: Data_out <= 16'h77C9	;
				14'b00110001010110: Data_out <= 16'h77CE	;
				14'b00110001010111: Data_out <= 16'h77D2	;
				14'b00110001011000: Data_out <= 16'h77D7	;
				14'b00110001011001: Data_out <= 16'h77DB	;
				14'b00110001011010: Data_out <= 16'h77E0	;
				14'b00110001011011: Data_out <= 16'h77E4	;
				14'b00110001011100: Data_out <= 16'h77E8	;
				14'b00110001011101: Data_out <= 16'h77ED	;
				14'b00110001011110: Data_out <= 16'h77F1	;
				14'b00110001011111: Data_out <= 16'h77F6	;
				14'b00110001100000: Data_out <= 16'h77FA	;
				14'b00110001100001: Data_out <= 16'h77FE	;
				14'b00110001100010: Data_out <= 16'h7803	;
				14'b00110001100011: Data_out <= 16'h7807	;
				14'b00110001100100: Data_out <= 16'h780B	;
				14'b00110001100101: Data_out <= 16'h7810	;
				14'b00110001100110: Data_out <= 16'h7814	;
				14'b00110001100111: Data_out <= 16'h7818	;
				14'b00110001101000: Data_out <= 16'h781D	;
				14'b00110001101001: Data_out <= 16'h7821	;
				14'b00110001101010: Data_out <= 16'h7825	;
				14'b00110001101011: Data_out <= 16'h782A	;
				14'b00110001101100: Data_out <= 16'h782E	;
				14'b00110001101101: Data_out <= 16'h7832	;
				14'b00110001101110: Data_out <= 16'h7837	;
				14'b00110001101111: Data_out <= 16'h783B	;
				14'b00110001110000: Data_out <= 16'h783F	;
				14'b00110001110001: Data_out <= 16'h7844	;
				14'b00110001110010: Data_out <= 16'h7848	;
				14'b00110001110011: Data_out <= 16'h784C	;
				14'b00110001110100: Data_out <= 16'h7851	;
				14'b00110001110101: Data_out <= 16'h7855	;
				14'b00110001110110: Data_out <= 16'h7859	;
				14'b00110001110111: Data_out <= 16'h785D	;
				14'b00110001111000: Data_out <= 16'h7862	;
				14'b00110001111001: Data_out <= 16'h7866	;
				14'b00110001111010: Data_out <= 16'h786A	;
				14'b00110001111011: Data_out <= 16'h786E	;
				14'b00110001111100: Data_out <= 16'h7873	;
				14'b00110001111101: Data_out <= 16'h7877	;
				14'b00110001111110: Data_out <= 16'h787B	;
				14'b00110001111111: Data_out <= 16'h787F	;
				14'b00110010000000: Data_out <= 16'h7884	;
				14'b00110010000001: Data_out <= 16'h7888	;
				14'b00110010000010: Data_out <= 16'h788C	;
				14'b00110010000011: Data_out <= 16'h7890	;
				14'b00110010000100: Data_out <= 16'h7895	;
				14'b00110010000101: Data_out <= 16'h7899	;
				14'b00110010000110: Data_out <= 16'h789D	;
				14'b00110010000111: Data_out <= 16'h78A1	;
				14'b00110010001000: Data_out <= 16'h78A5	;
				14'b00110010001001: Data_out <= 16'h78AA	;
				14'b00110010001010: Data_out <= 16'h78AE	;
				14'b00110010001011: Data_out <= 16'h78B2	;
				14'b00110010001100: Data_out <= 16'h78B6	;
				14'b00110010001101: Data_out <= 16'h78BA	;
				14'b00110010001110: Data_out <= 16'h78BE	;
				14'b00110010001111: Data_out <= 16'h78C3	;
				14'b00110010010000: Data_out <= 16'h78C7	;
				14'b00110010010001: Data_out <= 16'h78CB	;
				14'b00110010010010: Data_out <= 16'h78CF	;
				14'b00110010010011: Data_out <= 16'h78D3	;
				14'b00110010010100: Data_out <= 16'h78D7	;
				14'b00110010010101: Data_out <= 16'h78DC	;
				14'b00110010010110: Data_out <= 16'h78E0	;
				14'b00110010010111: Data_out <= 16'h78E4	;
				14'b00110010011000: Data_out <= 16'h78E8	;
				14'b00110010011001: Data_out <= 16'h78EC	;
				14'b00110010011010: Data_out <= 16'h78F0	;
				14'b00110010011011: Data_out <= 16'h78F4	;
				14'b00110010011100: Data_out <= 16'h78F8	;
				14'b00110010011101: Data_out <= 16'h78FD	;
				14'b00110010011110: Data_out <= 16'h7901	;
				14'b00110010011111: Data_out <= 16'h7905	;
				14'b00110010100000: Data_out <= 16'h7909	;
				14'b00110010100001: Data_out <= 16'h790D	;
				14'b00110010100010: Data_out <= 16'h7911	;
				14'b00110010100011: Data_out <= 16'h7915	;
				14'b00110010100100: Data_out <= 16'h7919	;
				14'b00110010100101: Data_out <= 16'h791D	;
				14'b00110010100110: Data_out <= 16'h7921	;
				14'b00110010100111: Data_out <= 16'h7925	;
				14'b00110010101000: Data_out <= 16'h7929	;
				14'b00110010101001: Data_out <= 16'h792D	;
				14'b00110010101010: Data_out <= 16'h7931	;
				14'b00110010101011: Data_out <= 16'h7936	;
				14'b00110010101100: Data_out <= 16'h793A	;
				14'b00110010101101: Data_out <= 16'h793E	;
				14'b00110010101110: Data_out <= 16'h7942	;
				14'b00110010101111: Data_out <= 16'h7946	;
				14'b00110010110000: Data_out <= 16'h794A	;
				14'b00110010110001: Data_out <= 16'h794E	;
				14'b00110010110010: Data_out <= 16'h7952	;
				14'b00110010110011: Data_out <= 16'h7956	;
				14'b00110010110100: Data_out <= 16'h795A	;
				14'b00110010110101: Data_out <= 16'h795E	;
				14'b00110010110110: Data_out <= 16'h7962	;
				14'b00110010110111: Data_out <= 16'h7966	;
				14'b00110010111000: Data_out <= 16'h796A	;
				14'b00110010111001: Data_out <= 16'h796E	;
				14'b00110010111010: Data_out <= 16'h7972	;
				14'b00110010111011: Data_out <= 16'h7976	;
				14'b00110010111100: Data_out <= 16'h7979	;
				14'b00110010111101: Data_out <= 16'h797D	;
				14'b00110010111110: Data_out <= 16'h7981	;
				14'b00110010111111: Data_out <= 16'h7985	;
				14'b00110011000000: Data_out <= 16'h7989	;
				14'b00110011000001: Data_out <= 16'h798D	;
				14'b00110011000010: Data_out <= 16'h7991	;
				14'b00110011000011: Data_out <= 16'h7995	;
				14'b00110011000100: Data_out <= 16'h7999	;
				14'b00110011000101: Data_out <= 16'h799D	;
				14'b00110011000110: Data_out <= 16'h79A1	;
				14'b00110011000111: Data_out <= 16'h79A5	;
				14'b00110011001000: Data_out <= 16'h79A9	;
				14'b00110011001001: Data_out <= 16'h79AD	;
				14'b00110011001010: Data_out <= 16'h79B0	;
				14'b00110011001011: Data_out <= 16'h79B4	;
				14'b00110011001100: Data_out <= 16'h79B8	;
				14'b00110011001101: Data_out <= 16'h79BC	;
				14'b00110011001110: Data_out <= 16'h79C0	;
				14'b00110011001111: Data_out <= 16'h79C4	;
				14'b00110011010000: Data_out <= 16'h79C8	;
				14'b00110011010001: Data_out <= 16'h79CC	;
				14'b00110011010010: Data_out <= 16'h79CF	;
				14'b00110011010011: Data_out <= 16'h79D3	;
				14'b00110011010100: Data_out <= 16'h79D7	;
				14'b00110011010101: Data_out <= 16'h79DB	;
				14'b00110011010110: Data_out <= 16'h79DF	;
				14'b00110011010111: Data_out <= 16'h79E3	;
				14'b00110011011000: Data_out <= 16'h79E7	;
				14'b00110011011001: Data_out <= 16'h79EA	;
				14'b00110011011010: Data_out <= 16'h79EE	;
				14'b00110011011011: Data_out <= 16'h79F2	;
				14'b00110011011100: Data_out <= 16'h79F6	;
				14'b00110011011101: Data_out <= 16'h79FA	;
				14'b00110011011110: Data_out <= 16'h79FD	;
				14'b00110011011111: Data_out <= 16'h7A01	;
				14'b00110011100000: Data_out <= 16'h7A05	;
				14'b00110011100001: Data_out <= 16'h7A09	;
				14'b00110011100010: Data_out <= 16'h7A0D	;
				14'b00110011100011: Data_out <= 16'h7A10	;
				14'b00110011100100: Data_out <= 16'h7A14	;
				14'b00110011100101: Data_out <= 16'h7A18	;
				14'b00110011100110: Data_out <= 16'h7A1C	;
				14'b00110011100111: Data_out <= 16'h7A20	;
				14'b00110011101000: Data_out <= 16'h7A23	;
				14'b00110011101001: Data_out <= 16'h7A27	;
				14'b00110011101010: Data_out <= 16'h7A2B	;
				14'b00110011101011: Data_out <= 16'h7A2F	;
				14'b00110011101100: Data_out <= 16'h7A32	;
				14'b00110011101101: Data_out <= 16'h7A36	;
				14'b00110011101110: Data_out <= 16'h7A3A	;
				14'b00110011101111: Data_out <= 16'h7A3D	;
				14'b00110011110000: Data_out <= 16'h7A41	;
				14'b00110011110001: Data_out <= 16'h7A45	;
				14'b00110011110010: Data_out <= 16'h7A49	;
				14'b00110011110011: Data_out <= 16'h7A4C	;
				14'b00110011110100: Data_out <= 16'h7A50	;
				14'b00110011110101: Data_out <= 16'h7A54	;
				14'b00110011110110: Data_out <= 16'h7A57	;
				14'b00110011110111: Data_out <= 16'h7A5B	;
				14'b00110011111000: Data_out <= 16'h7A5F	;
				14'b00110011111001: Data_out <= 16'h7A63	;
				14'b00110011111010: Data_out <= 16'h7A66	;
				14'b00110011111011: Data_out <= 16'h7A6A	;
				14'b00110011111100: Data_out <= 16'h7A6E	;
				14'b00110011111101: Data_out <= 16'h7A71	;
				14'b00110011111110: Data_out <= 16'h7A75	;
				14'b00110011111111: Data_out <= 16'h7A79	;
				14'b00110100000000: Data_out <= 16'h7A7C	;
				14'b00110100000001: Data_out <= 16'h7A80	;
				14'b00110100000010: Data_out <= 16'h7A83	;
				14'b00110100000011: Data_out <= 16'h7A87	;
				14'b00110100000100: Data_out <= 16'h7A8B	;
				14'b00110100000101: Data_out <= 16'h7A8E	;
				14'b00110100000110: Data_out <= 16'h7A92	;
				14'b00110100000111: Data_out <= 16'h7A96	;
				14'b00110100001000: Data_out <= 16'h7A99	;
				14'b00110100001001: Data_out <= 16'h7A9D	;
				14'b00110100001010: Data_out <= 16'h7AA0	;
				14'b00110100001011: Data_out <= 16'h7AA4	;
				14'b00110100001100: Data_out <= 16'h7AA8	;
				14'b00110100001101: Data_out <= 16'h7AAB	;
				14'b00110100001110: Data_out <= 16'h7AAF	;
				14'b00110100001111: Data_out <= 16'h7AB2	;
				14'b00110100010000: Data_out <= 16'h7AB6	;
				14'b00110100010001: Data_out <= 16'h7ABA	;
				14'b00110100010010: Data_out <= 16'h7ABD	;
				14'b00110100010011: Data_out <= 16'h7AC1	;
				14'b00110100010100: Data_out <= 16'h7AC4	;
				14'b00110100010101: Data_out <= 16'h7AC8	;
				14'b00110100010110: Data_out <= 16'h7ACB	;
				14'b00110100010111: Data_out <= 16'h7ACF	;
				14'b00110100011000: Data_out <= 16'h7AD2	;
				14'b00110100011001: Data_out <= 16'h7AD6	;
				14'b00110100011010: Data_out <= 16'h7AD9	;
				14'b00110100011011: Data_out <= 16'h7ADD	;
				14'b00110100011100: Data_out <= 16'h7AE0	;
				14'b00110100011101: Data_out <= 16'h7AE4	;
				14'b00110100011110: Data_out <= 16'h7AE8	;
				14'b00110100011111: Data_out <= 16'h7AEB	;
				14'b00110100100000: Data_out <= 16'h7AEF	;
				14'b00110100100001: Data_out <= 16'h7AF2	;
				14'b00110100100010: Data_out <= 16'h7AF6	;
				14'b00110100100011: Data_out <= 16'h7AF9	;
				14'b00110100100100: Data_out <= 16'h7AFC	;
				14'b00110100100101: Data_out <= 16'h7B00	;
				14'b00110100100110: Data_out <= 16'h7B03	;
				14'b00110100100111: Data_out <= 16'h7B07	;
				14'b00110100101000: Data_out <= 16'h7B0A	;
				14'b00110100101001: Data_out <= 16'h7B0E	;
				14'b00110100101010: Data_out <= 16'h7B11	;
				14'b00110100101011: Data_out <= 16'h7B15	;
				14'b00110100101100: Data_out <= 16'h7B18	;
				14'b00110100101101: Data_out <= 16'h7B1C	;
				14'b00110100101110: Data_out <= 16'h7B1F	;
				14'b00110100101111: Data_out <= 16'h7B23	;
				14'b00110100110000: Data_out <= 16'h7B26	;
				14'b00110100110001: Data_out <= 16'h7B29	;
				14'b00110100110010: Data_out <= 16'h7B2D	;
				14'b00110100110011: Data_out <= 16'h7B30	;
				14'b00110100110100: Data_out <= 16'h7B34	;
				14'b00110100110101: Data_out <= 16'h7B37	;
				14'b00110100110110: Data_out <= 16'h7B3A	;
				14'b00110100110111: Data_out <= 16'h7B3E	;
				14'b00110100111000: Data_out <= 16'h7B41	;
				14'b00110100111001: Data_out <= 16'h7B45	;
				14'b00110100111010: Data_out <= 16'h7B48	;
				14'b00110100111011: Data_out <= 16'h7B4B	;
				14'b00110100111100: Data_out <= 16'h7B4F	;
				14'b00110100111101: Data_out <= 16'h7B52	;
				14'b00110100111110: Data_out <= 16'h7B55	;
				14'b00110100111111: Data_out <= 16'h7B59	;
				14'b00110101000000: Data_out <= 16'h7B5C	;
				14'b00110101000001: Data_out <= 16'h7B5F	;
				14'b00110101000010: Data_out <= 16'h7B63	;
				14'b00110101000011: Data_out <= 16'h7B66	;
				14'b00110101000100: Data_out <= 16'h7B6A	;
				14'b00110101000101: Data_out <= 16'h7B6D	;
				14'b00110101000110: Data_out <= 16'h7B70	;
				14'b00110101000111: Data_out <= 16'h7B73	;
				14'b00110101001000: Data_out <= 16'h7B77	;
				14'b00110101001001: Data_out <= 16'h7B7A	;
				14'b00110101001010: Data_out <= 16'h7B7D	;
				14'b00110101001011: Data_out <= 16'h7B81	;
				14'b00110101001100: Data_out <= 16'h7B84	;
				14'b00110101001101: Data_out <= 16'h7B87	;
				14'b00110101001110: Data_out <= 16'h7B8B	;
				14'b00110101001111: Data_out <= 16'h7B8E	;
				14'b00110101010000: Data_out <= 16'h7B91	;
				14'b00110101010001: Data_out <= 16'h7B94	;
				14'b00110101010010: Data_out <= 16'h7B98	;
				14'b00110101010011: Data_out <= 16'h7B9B	;
				14'b00110101010100: Data_out <= 16'h7B9E	;
				14'b00110101010101: Data_out <= 16'h7BA2	;
				14'b00110101010110: Data_out <= 16'h7BA5	;
				14'b00110101010111: Data_out <= 16'h7BA8	;
				14'b00110101011000: Data_out <= 16'h7BAB	;
				14'b00110101011001: Data_out <= 16'h7BAE	;
				14'b00110101011010: Data_out <= 16'h7BB2	;
				14'b00110101011011: Data_out <= 16'h7BB5	;
				14'b00110101011100: Data_out <= 16'h7BB8	;
				14'b00110101011101: Data_out <= 16'h7BBB	;
				14'b00110101011110: Data_out <= 16'h7BBF	;
				14'b00110101011111: Data_out <= 16'h7BC2	;
				14'b00110101100000: Data_out <= 16'h7BC5	;
				14'b00110101100001: Data_out <= 16'h7BC8	;
				14'b00110101100010: Data_out <= 16'h7BCB	;
				14'b00110101100011: Data_out <= 16'h7BCF	;
				14'b00110101100100: Data_out <= 16'h7BD2	;
				14'b00110101100101: Data_out <= 16'h7BD5	;
				14'b00110101100110: Data_out <= 16'h7BD8	;
				14'b00110101100111: Data_out <= 16'h7BDB	;
				14'b00110101101000: Data_out <= 16'h7BDE	;
				14'b00110101101001: Data_out <= 16'h7BE2	;
				14'b00110101101010: Data_out <= 16'h7BE5	;
				14'b00110101101011: Data_out <= 16'h7BE8	;
				14'b00110101101100: Data_out <= 16'h7BEB	;
				14'b00110101101101: Data_out <= 16'h7BEE	;
				14'b00110101101110: Data_out <= 16'h7BF1	;
				14'b00110101101111: Data_out <= 16'h7BF5	;
				14'b00110101110000: Data_out <= 16'h7BF8	;
				14'b00110101110001: Data_out <= 16'h7BFB	;
				14'b00110101110010: Data_out <= 16'h7BFE	;
				14'b00110101110011: Data_out <= 16'h7C01	;
				14'b00110101110100: Data_out <= 16'h7C04	;
				14'b00110101110101: Data_out <= 16'h7C07	;
				14'b00110101110110: Data_out <= 16'h7C0A	;
				14'b00110101110111: Data_out <= 16'h7C0D	;
				14'b00110101111000: Data_out <= 16'h7C11	;
				14'b00110101111001: Data_out <= 16'h7C14	;
				14'b00110101111010: Data_out <= 16'h7C17	;
				14'b00110101111011: Data_out <= 16'h7C1A	;
				14'b00110101111100: Data_out <= 16'h7C1D	;
				14'b00110101111101: Data_out <= 16'h7C20	;
				14'b00110101111110: Data_out <= 16'h7C23	;
				14'b00110101111111: Data_out <= 16'h7C26	;
				14'b00110110000000: Data_out <= 16'h7C29	;
				14'b00110110000001: Data_out <= 16'h7C2C	;
				14'b00110110000010: Data_out <= 16'h7C2F	;
				14'b00110110000011: Data_out <= 16'h7C32	;
				14'b00110110000100: Data_out <= 16'h7C35	;
				14'b00110110000101: Data_out <= 16'h7C38	;
				14'b00110110000110: Data_out <= 16'h7C3B	;
				14'b00110110000111: Data_out <= 16'h7C3E	;
				14'b00110110001000: Data_out <= 16'h7C41	;
				14'b00110110001001: Data_out <= 16'h7C44	;
				14'b00110110001010: Data_out <= 16'h7C47	;
				14'b00110110001011: Data_out <= 16'h7C4A	;
				14'b00110110001100: Data_out <= 16'h7C4D	;
				14'b00110110001101: Data_out <= 16'h7C50	;
				14'b00110110001110: Data_out <= 16'h7C53	;
				14'b00110110001111: Data_out <= 16'h7C56	;
				14'b00110110010000: Data_out <= 16'h7C59	;
				14'b00110110010001: Data_out <= 16'h7C5C	;
				14'b00110110010010: Data_out <= 16'h7C5F	;
				14'b00110110010011: Data_out <= 16'h7C62	;
				14'b00110110010100: Data_out <= 16'h7C65	;
				14'b00110110010101: Data_out <= 16'h7C68	;
				14'b00110110010110: Data_out <= 16'h7C6B	;
				14'b00110110010111: Data_out <= 16'h7C6E	;
				14'b00110110011000: Data_out <= 16'h7C71	;
				14'b00110110011001: Data_out <= 16'h7C74	;
				14'b00110110011010: Data_out <= 16'h7C77	;
				14'b00110110011011: Data_out <= 16'h7C7A	;
				14'b00110110011100: Data_out <= 16'h7C7D	;
				14'b00110110011101: Data_out <= 16'h7C80	;
				14'b00110110011110: Data_out <= 16'h7C83	;
				14'b00110110011111: Data_out <= 16'h7C86	;
				14'b00110110100000: Data_out <= 16'h7C88	;
				14'b00110110100001: Data_out <= 16'h7C8B	;
				14'b00110110100010: Data_out <= 16'h7C8E	;
				14'b00110110100011: Data_out <= 16'h7C91	;
				14'b00110110100100: Data_out <= 16'h7C94	;
				14'b00110110100101: Data_out <= 16'h7C97	;
				14'b00110110100110: Data_out <= 16'h7C9A	;
				14'b00110110100111: Data_out <= 16'h7C9D	;
				14'b00110110101000: Data_out <= 16'h7CA0	;
				14'b00110110101001: Data_out <= 16'h7CA2	;
				14'b00110110101010: Data_out <= 16'h7CA5	;
				14'b00110110101011: Data_out <= 16'h7CA8	;
				14'b00110110101100: Data_out <= 16'h7CAB	;
				14'b00110110101101: Data_out <= 16'h7CAE	;
				14'b00110110101110: Data_out <= 16'h7CB1	;
				14'b00110110101111: Data_out <= 16'h7CB3	;
				14'b00110110110000: Data_out <= 16'h7CB6	;
				14'b00110110110001: Data_out <= 16'h7CB9	;
				14'b00110110110010: Data_out <= 16'h7CBC	;
				14'b00110110110011: Data_out <= 16'h7CBF	;
				14'b00110110110100: Data_out <= 16'h7CC2	;
				14'b00110110110101: Data_out <= 16'h7CC4	;
				14'b00110110110110: Data_out <= 16'h7CC7	;
				14'b00110110110111: Data_out <= 16'h7CCA	;
				14'b00110110111000: Data_out <= 16'h7CCD	;
				14'b00110110111001: Data_out <= 16'h7CD0	;
				14'b00110110111010: Data_out <= 16'h7CD2	;
				14'b00110110111011: Data_out <= 16'h7CD5	;
				14'b00110110111100: Data_out <= 16'h7CD8	;
				14'b00110110111101: Data_out <= 16'h7CDB	;
				14'b00110110111110: Data_out <= 16'h7CDD	;
				14'b00110110111111: Data_out <= 16'h7CE0	;
				14'b00110111000000: Data_out <= 16'h7CE3	;
				14'b00110111000001: Data_out <= 16'h7CE6	;
				14'b00110111000010: Data_out <= 16'h7CE8	;
				14'b00110111000011: Data_out <= 16'h7CEB	;
				14'b00110111000100: Data_out <= 16'h7CEE	;
				14'b00110111000101: Data_out <= 16'h7CF1	;
				14'b00110111000110: Data_out <= 16'h7CF3	;
				14'b00110111000111: Data_out <= 16'h7CF6	;
				14'b00110111001000: Data_out <= 16'h7CF9	;
				14'b00110111001001: Data_out <= 16'h7CFC	;
				14'b00110111001010: Data_out <= 16'h7CFE	;
				14'b00110111001011: Data_out <= 16'h7D01	;
				14'b00110111001100: Data_out <= 16'h7D04	;
				14'b00110111001101: Data_out <= 16'h7D06	;
				14'b00110111001110: Data_out <= 16'h7D09	;
				14'b00110111001111: Data_out <= 16'h7D0C	;
				14'b00110111010000: Data_out <= 16'h7D0E	;
				14'b00110111010001: Data_out <= 16'h7D11	;
				14'b00110111010010: Data_out <= 16'h7D14	;
				14'b00110111010011: Data_out <= 16'h7D16	;
				14'b00110111010100: Data_out <= 16'h7D19	;
				14'b00110111010101: Data_out <= 16'h7D1C	;
				14'b00110111010110: Data_out <= 16'h7D1E	;
				14'b00110111010111: Data_out <= 16'h7D21	;
				14'b00110111011000: Data_out <= 16'h7D24	;
				14'b00110111011001: Data_out <= 16'h7D26	;
				14'b00110111011010: Data_out <= 16'h7D29	;
				14'b00110111011011: Data_out <= 16'h7D2C	;
				14'b00110111011100: Data_out <= 16'h7D2E	;
				14'b00110111011101: Data_out <= 16'h7D31	;
				14'b00110111011110: Data_out <= 16'h7D33	;
				14'b00110111011111: Data_out <= 16'h7D36	;
				14'b00110111100000: Data_out <= 16'h7D39	;
				14'b00110111100001: Data_out <= 16'h7D3B	;
				14'b00110111100010: Data_out <= 16'h7D3E	;
				14'b00110111100011: Data_out <= 16'h7D40	;
				14'b00110111100100: Data_out <= 16'h7D43	;
				14'b00110111100101: Data_out <= 16'h7D46	;
				14'b00110111100110: Data_out <= 16'h7D48	;
				14'b00110111100111: Data_out <= 16'h7D4B	;
				14'b00110111101000: Data_out <= 16'h7D4D	;
				14'b00110111101001: Data_out <= 16'h7D50	;
				14'b00110111101010: Data_out <= 16'h7D52	;
				14'b00110111101011: Data_out <= 16'h7D55	;
				14'b00110111101100: Data_out <= 16'h7D58	;
				14'b00110111101101: Data_out <= 16'h7D5A	;
				14'b00110111101110: Data_out <= 16'h7D5D	;
				14'b00110111101111: Data_out <= 16'h7D5F	;
				14'b00110111110000: Data_out <= 16'h7D62	;
				14'b00110111110001: Data_out <= 16'h7D64	;
				14'b00110111110010: Data_out <= 16'h7D67	;
				14'b00110111110011: Data_out <= 16'h7D69	;
				14'b00110111110100: Data_out <= 16'h7D6C	;
				14'b00110111110101: Data_out <= 16'h7D6E	;
				14'b00110111110110: Data_out <= 16'h7D71	;
				14'b00110111110111: Data_out <= 16'h7D73	;
				14'b00110111111000: Data_out <= 16'h7D76	;
				14'b00110111111001: Data_out <= 16'h7D78	;
				14'b00110111111010: Data_out <= 16'h7D7B	;
				14'b00110111111011: Data_out <= 16'h7D7D	;
				14'b00110111111100: Data_out <= 16'h7D80	;
				14'b00110111111101: Data_out <= 16'h7D82	;
				14'b00110111111110: Data_out <= 16'h7D85	;
				14'b00110111111111: Data_out <= 16'h7D87	;
				14'b00111000000000: Data_out <= 16'h7D89	;
				14'b00111000000001: Data_out <= 16'h7D8C	;
				14'b00111000000010: Data_out <= 16'h7D8E	;
				14'b00111000000011: Data_out <= 16'h7D91	;
				14'b00111000000100: Data_out <= 16'h7D93	;
				14'b00111000000101: Data_out <= 16'h7D96	;
				14'b00111000000110: Data_out <= 16'h7D98	;
				14'b00111000000111: Data_out <= 16'h7D9B	;
				14'b00111000001000: Data_out <= 16'h7D9D	;
				14'b00111000001001: Data_out <= 16'h7D9F	;
				14'b00111000001010: Data_out <= 16'h7DA2	;
				14'b00111000001011: Data_out <= 16'h7DA4	;
				14'b00111000001100: Data_out <= 16'h7DA7	;
				14'b00111000001101: Data_out <= 16'h7DA9	;
				14'b00111000001110: Data_out <= 16'h7DAB	;
				14'b00111000001111: Data_out <= 16'h7DAE	;
				14'b00111000010000: Data_out <= 16'h7DB0	;
				14'b00111000010001: Data_out <= 16'h7DB2	;
				14'b00111000010010: Data_out <= 16'h7DB5	;
				14'b00111000010011: Data_out <= 16'h7DB7	;
				14'b00111000010100: Data_out <= 16'h7DBA	;
				14'b00111000010101: Data_out <= 16'h7DBC	;
				14'b00111000010110: Data_out <= 16'h7DBE	;
				14'b00111000010111: Data_out <= 16'h7DC1	;
				14'b00111000011000: Data_out <= 16'h7DC3	;
				14'b00111000011001: Data_out <= 16'h7DC5	;
				14'b00111000011010: Data_out <= 16'h7DC8	;
				14'b00111000011011: Data_out <= 16'h7DCA	;
				14'b00111000011100: Data_out <= 16'h7DCC	;
				14'b00111000011101: Data_out <= 16'h7DCF	;
				14'b00111000011110: Data_out <= 16'h7DD1	;
				14'b00111000011111: Data_out <= 16'h7DD3	;
				14'b00111000100000: Data_out <= 16'h7DD6	;
				14'b00111000100001: Data_out <= 16'h7DD8	;
				14'b00111000100010: Data_out <= 16'h7DDA	;
				14'b00111000100011: Data_out <= 16'h7DDC	;
				14'b00111000100100: Data_out <= 16'h7DDF	;
				14'b00111000100101: Data_out <= 16'h7DE1	;
				14'b00111000100110: Data_out <= 16'h7DE3	;
				14'b00111000100111: Data_out <= 16'h7DE6	;
				14'b00111000101000: Data_out <= 16'h7DE8	;
				14'b00111000101001: Data_out <= 16'h7DEA	;
				14'b00111000101010: Data_out <= 16'h7DEC	;
				14'b00111000101011: Data_out <= 16'h7DEF	;
				14'b00111000101100: Data_out <= 16'h7DF1	;
				14'b00111000101101: Data_out <= 16'h7DF3	;
				14'b00111000101110: Data_out <= 16'h7DF5	;
				14'b00111000101111: Data_out <= 16'h7DF7	;
				14'b00111000110000: Data_out <= 16'h7DFA	;
				14'b00111000110001: Data_out <= 16'h7DFC	;
				14'b00111000110010: Data_out <= 16'h7DFE	;
				14'b00111000110011: Data_out <= 16'h7E00	;
				14'b00111000110100: Data_out <= 16'h7E03	;
				14'b00111000110101: Data_out <= 16'h7E05	;
				14'b00111000110110: Data_out <= 16'h7E07	;
				14'b00111000110111: Data_out <= 16'h7E09	;
				14'b00111000111000: Data_out <= 16'h7E0B	;
				14'b00111000111001: Data_out <= 16'h7E0E	;
				14'b00111000111010: Data_out <= 16'h7E10	;
				14'b00111000111011: Data_out <= 16'h7E12	;
				14'b00111000111100: Data_out <= 16'h7E14	;
				14'b00111000111101: Data_out <= 16'h7E16	;
				14'b00111000111110: Data_out <= 16'h7E18	;
				14'b00111000111111: Data_out <= 16'h7E1B	;
				14'b00111001000000: Data_out <= 16'h7E1D	;
				14'b00111001000001: Data_out <= 16'h7E1F	;
				14'b00111001000010: Data_out <= 16'h7E21	;
				14'b00111001000011: Data_out <= 16'h7E23	;
				14'b00111001000100: Data_out <= 16'h7E25	;
				14'b00111001000101: Data_out <= 16'h7E27	;
				14'b00111001000110: Data_out <= 16'h7E29	;
				14'b00111001000111: Data_out <= 16'h7E2C	;
				14'b00111001001000: Data_out <= 16'h7E2E	;
				14'b00111001001001: Data_out <= 16'h7E30	;
				14'b00111001001010: Data_out <= 16'h7E32	;
				14'b00111001001011: Data_out <= 16'h7E34	;
				14'b00111001001100: Data_out <= 16'h7E36	;
				14'b00111001001101: Data_out <= 16'h7E38	;
				14'b00111001001110: Data_out <= 16'h7E3A	;
				14'b00111001001111: Data_out <= 16'h7E3C	;
				14'b00111001010000: Data_out <= 16'h7E3E	;
				14'b00111001010001: Data_out <= 16'h7E41	;
				14'b00111001010010: Data_out <= 16'h7E43	;
				14'b00111001010011: Data_out <= 16'h7E45	;
				14'b00111001010100: Data_out <= 16'h7E47	;
				14'b00111001010101: Data_out <= 16'h7E49	;
				14'b00111001010110: Data_out <= 16'h7E4B	;
				14'b00111001010111: Data_out <= 16'h7E4D	;
				14'b00111001011000: Data_out <= 16'h7E4F	;
				14'b00111001011001: Data_out <= 16'h7E51	;
				14'b00111001011010: Data_out <= 16'h7E53	;
				14'b00111001011011: Data_out <= 16'h7E55	;
				14'b00111001011100: Data_out <= 16'h7E57	;
				14'b00111001011101: Data_out <= 16'h7E59	;
				14'b00111001011110: Data_out <= 16'h7E5B	;
				14'b00111001011111: Data_out <= 16'h7E5D	;
				14'b00111001100000: Data_out <= 16'h7E5F	;
				14'b00111001100001: Data_out <= 16'h7E61	;
				14'b00111001100010: Data_out <= 16'h7E63	;
				14'b00111001100011: Data_out <= 16'h7E65	;
				14'b00111001100100: Data_out <= 16'h7E67	;
				14'b00111001100101: Data_out <= 16'h7E69	;
				14'b00111001100110: Data_out <= 16'h7E6B	;
				14'b00111001100111: Data_out <= 16'h7E6D	;
				14'b00111001101000: Data_out <= 16'h7E6F	;
				14'b00111001101001: Data_out <= 16'h7E71	;
				14'b00111001101010: Data_out <= 16'h7E73	;
				14'b00111001101011: Data_out <= 16'h7E75	;
				14'b00111001101100: Data_out <= 16'h7E77	;
				14'b00111001101101: Data_out <= 16'h7E79	;
				14'b00111001101110: Data_out <= 16'h7E7A	;
				14'b00111001101111: Data_out <= 16'h7E7C	;
				14'b00111001110000: Data_out <= 16'h7E7E	;
				14'b00111001110001: Data_out <= 16'h7E80	;
				14'b00111001110010: Data_out <= 16'h7E82	;
				14'b00111001110011: Data_out <= 16'h7E84	;
				14'b00111001110100: Data_out <= 16'h7E86	;
				14'b00111001110101: Data_out <= 16'h7E88	;
				14'b00111001110110: Data_out <= 16'h7E8A	;
				14'b00111001110111: Data_out <= 16'h7E8C	;
				14'b00111001111000: Data_out <= 16'h7E8E	;
				14'b00111001111001: Data_out <= 16'h7E8F	;
				14'b00111001111010: Data_out <= 16'h7E91	;
				14'b00111001111011: Data_out <= 16'h7E93	;
				14'b00111001111100: Data_out <= 16'h7E95	;
				14'b00111001111101: Data_out <= 16'h7E97	;
				14'b00111001111110: Data_out <= 16'h7E99	;
				14'b00111001111111: Data_out <= 16'h7E9B	;
				14'b00111010000000: Data_out <= 16'h7E9C	;
				14'b00111010000001: Data_out <= 16'h7E9E	;
				14'b00111010000010: Data_out <= 16'h7EA0	;
				14'b00111010000011: Data_out <= 16'h7EA2	;
				14'b00111010000100: Data_out <= 16'h7EA4	;
				14'b00111010000101: Data_out <= 16'h7EA6	;
				14'b00111010000110: Data_out <= 16'h7EA7	;
				14'b00111010000111: Data_out <= 16'h7EA9	;
				14'b00111010001000: Data_out <= 16'h7EAB	;
				14'b00111010001001: Data_out <= 16'h7EAD	;
				14'b00111010001010: Data_out <= 16'h7EAF	;
				14'b00111010001011: Data_out <= 16'h7EB0	;
				14'b00111010001100: Data_out <= 16'h7EB2	;
				14'b00111010001101: Data_out <= 16'h7EB4	;
				14'b00111010001110: Data_out <= 16'h7EB6	;
				14'b00111010001111: Data_out <= 16'h7EB8	;
				14'b00111010010000: Data_out <= 16'h7EB9	;
				14'b00111010010001: Data_out <= 16'h7EBB	;
				14'b00111010010010: Data_out <= 16'h7EBD	;
				14'b00111010010011: Data_out <= 16'h7EBF	;
				14'b00111010010100: Data_out <= 16'h7EC0	;
				14'b00111010010101: Data_out <= 16'h7EC2	;
				14'b00111010010110: Data_out <= 16'h7EC4	;
				14'b00111010010111: Data_out <= 16'h7EC6	;
				14'b00111010011000: Data_out <= 16'h7EC7	;
				14'b00111010011001: Data_out <= 16'h7EC9	;
				14'b00111010011010: Data_out <= 16'h7ECB	;
				14'b00111010011011: Data_out <= 16'h7ECC	;
				14'b00111010011100: Data_out <= 16'h7ECE	;
				14'b00111010011101: Data_out <= 16'h7ED0	;
				14'b00111010011110: Data_out <= 16'h7ED2	;
				14'b00111010011111: Data_out <= 16'h7ED3	;
				14'b00111010100000: Data_out <= 16'h7ED5	;
				14'b00111010100001: Data_out <= 16'h7ED7	;
				14'b00111010100010: Data_out <= 16'h7ED8	;
				14'b00111010100011: Data_out <= 16'h7EDA	;
				14'b00111010100100: Data_out <= 16'h7EDC	;
				14'b00111010100101: Data_out <= 16'h7EDD	;
				14'b00111010100110: Data_out <= 16'h7EDF	;
				14'b00111010100111: Data_out <= 16'h7EE1	;
				14'b00111010101000: Data_out <= 16'h7EE2	;
				14'b00111010101001: Data_out <= 16'h7EE4	;
				14'b00111010101010: Data_out <= 16'h7EE6	;
				14'b00111010101011: Data_out <= 16'h7EE7	;
				14'b00111010101100: Data_out <= 16'h7EE9	;
				14'b00111010101101: Data_out <= 16'h7EEB	;
				14'b00111010101110: Data_out <= 16'h7EEC	;
				14'b00111010101111: Data_out <= 16'h7EEE	;
				14'b00111010110000: Data_out <= 16'h7EEF	;
				14'b00111010110001: Data_out <= 16'h7EF1	;
				14'b00111010110010: Data_out <= 16'h7EF3	;
				14'b00111010110011: Data_out <= 16'h7EF4	;
				14'b00111010110100: Data_out <= 16'h7EF6	;
				14'b00111010110101: Data_out <= 16'h7EF7	;
				14'b00111010110110: Data_out <= 16'h7EF9	;
				14'b00111010110111: Data_out <= 16'h7EFB	;
				14'b00111010111000: Data_out <= 16'h7EFC	;
				14'b00111010111001: Data_out <= 16'h7EFE	;
				14'b00111010111010: Data_out <= 16'h7EFF	;
				14'b00111010111011: Data_out <= 16'h7F01	;
				14'b00111010111100: Data_out <= 16'h7F02	;
				14'b00111010111101: Data_out <= 16'h7F04	;
				14'b00111010111110: Data_out <= 16'h7F06	;
				14'b00111010111111: Data_out <= 16'h7F07	;
				14'b00111011000000: Data_out <= 16'h7F09	;
				14'b00111011000001: Data_out <= 16'h7F0A	;
				14'b00111011000010: Data_out <= 16'h7F0C	;
				14'b00111011000011: Data_out <= 16'h7F0D	;
				14'b00111011000100: Data_out <= 16'h7F0F	;
				14'b00111011000101: Data_out <= 16'h7F10	;
				14'b00111011000110: Data_out <= 16'h7F12	;
				14'b00111011000111: Data_out <= 16'h7F13	;
				14'b00111011001000: Data_out <= 16'h7F15	;
				14'b00111011001001: Data_out <= 16'h7F16	;
				14'b00111011001010: Data_out <= 16'h7F18	;
				14'b00111011001011: Data_out <= 16'h7F19	;
				14'b00111011001100: Data_out <= 16'h7F1B	;
				14'b00111011001101: Data_out <= 16'h7F1C	;
				14'b00111011001110: Data_out <= 16'h7F1E	;
				14'b00111011001111: Data_out <= 16'h7F1F	;
				14'b00111011010000: Data_out <= 16'h7F21	;
				14'b00111011010001: Data_out <= 16'h7F22	;
				14'b00111011010010: Data_out <= 16'h7F24	;
				14'b00111011010011: Data_out <= 16'h7F25	;
				14'b00111011010100: Data_out <= 16'h7F26	;
				14'b00111011010101: Data_out <= 16'h7F28	;
				14'b00111011010110: Data_out <= 16'h7F29	;
				14'b00111011010111: Data_out <= 16'h7F2B	;
				14'b00111011011000: Data_out <= 16'h7F2C	;
				14'b00111011011001: Data_out <= 16'h7F2E	;
				14'b00111011011010: Data_out <= 16'h7F2F	;
				14'b00111011011011: Data_out <= 16'h7F30	;
				14'b00111011011100: Data_out <= 16'h7F32	;
				14'b00111011011101: Data_out <= 16'h7F33	;
				14'b00111011011110: Data_out <= 16'h7F35	;
				14'b00111011011111: Data_out <= 16'h7F36	;
				14'b00111011100000: Data_out <= 16'h7F37	;
				14'b00111011100001: Data_out <= 16'h7F39	;
				14'b00111011100010: Data_out <= 16'h7F3A	;
				14'b00111011100011: Data_out <= 16'h7F3C	;
				14'b00111011100100: Data_out <= 16'h7F3D	;
				14'b00111011100101: Data_out <= 16'h7F3E	;
				14'b00111011100110: Data_out <= 16'h7F40	;
				14'b00111011100111: Data_out <= 16'h7F41	;
				14'b00111011101000: Data_out <= 16'h7F42	;
				14'b00111011101001: Data_out <= 16'h7F44	;
				14'b00111011101010: Data_out <= 16'h7F45	;
				14'b00111011101011: Data_out <= 16'h7F46	;
				14'b00111011101100: Data_out <= 16'h7F48	;
				14'b00111011101101: Data_out <= 16'h7F49	;
				14'b00111011101110: Data_out <= 16'h7F4A	;
				14'b00111011101111: Data_out <= 16'h7F4C	;
				14'b00111011110000: Data_out <= 16'h7F4D	;
				14'b00111011110001: Data_out <= 16'h7F4E	;
				14'b00111011110010: Data_out <= 16'h7F50	;
				14'b00111011110011: Data_out <= 16'h7F51	;
				14'b00111011110100: Data_out <= 16'h7F52	;
				14'b00111011110101: Data_out <= 16'h7F53	;
				14'b00111011110110: Data_out <= 16'h7F55	;
				14'b00111011110111: Data_out <= 16'h7F56	;
				14'b00111011111000: Data_out <= 16'h7F57	;
				14'b00111011111001: Data_out <= 16'h7F59	;
				14'b00111011111010: Data_out <= 16'h7F5A	;
				14'b00111011111011: Data_out <= 16'h7F5B	;
				14'b00111011111100: Data_out <= 16'h7F5C	;
				14'b00111011111101: Data_out <= 16'h7F5E	;
				14'b00111011111110: Data_out <= 16'h7F5F	;
				14'b00111011111111: Data_out <= 16'h7F60	;
				14'b00111100000000: Data_out <= 16'h7F61	;
				14'b00111100000001: Data_out <= 16'h7F63	;
				14'b00111100000010: Data_out <= 16'h7F64	;
				14'b00111100000011: Data_out <= 16'h7F65	;
				14'b00111100000100: Data_out <= 16'h7F66	;
				14'b00111100000101: Data_out <= 16'h7F67	;
				14'b00111100000110: Data_out <= 16'h7F69	;
				14'b00111100000111: Data_out <= 16'h7F6A	;
				14'b00111100001000: Data_out <= 16'h7F6B	;
				14'b00111100001001: Data_out <= 16'h7F6C	;
				14'b00111100001010: Data_out <= 16'h7F6D	;
				14'b00111100001011: Data_out <= 16'h7F6F	;
				14'b00111100001100: Data_out <= 16'h7F70	;
				14'b00111100001101: Data_out <= 16'h7F71	;
				14'b00111100001110: Data_out <= 16'h7F72	;
				14'b00111100001111: Data_out <= 16'h7F73	;
				14'b00111100010000: Data_out <= 16'h7F74	;
				14'b00111100010001: Data_out <= 16'h7F76	;
				14'b00111100010010: Data_out <= 16'h7F77	;
				14'b00111100010011: Data_out <= 16'h7F78	;
				14'b00111100010100: Data_out <= 16'h7F79	;
				14'b00111100010101: Data_out <= 16'h7F7A	;
				14'b00111100010110: Data_out <= 16'h7F7B	;
				14'b00111100010111: Data_out <= 16'h7F7C	;
				14'b00111100011000: Data_out <= 16'h7F7D	;
				14'b00111100011001: Data_out <= 16'h7F7F	;
				14'b00111100011010: Data_out <= 16'h7F80	;
				14'b00111100011011: Data_out <= 16'h7F81	;
				14'b00111100011100: Data_out <= 16'h7F82	;
				14'b00111100011101: Data_out <= 16'h7F83	;
				14'b00111100011110: Data_out <= 16'h7F84	;
				14'b00111100011111: Data_out <= 16'h7F85	;
				14'b00111100100000: Data_out <= 16'h7F86	;
				14'b00111100100001: Data_out <= 16'h7F87	;
				14'b00111100100010: Data_out <= 16'h7F88	;
				14'b00111100100011: Data_out <= 16'h7F89	;
				14'b00111100100100: Data_out <= 16'h7F8B	;
				14'b00111100100101: Data_out <= 16'h7F8C	;
				14'b00111100100110: Data_out <= 16'h7F8D	;
				14'b00111100100111: Data_out <= 16'h7F8E	;
				14'b00111100101000: Data_out <= 16'h7F8F	;
				14'b00111100101001: Data_out <= 16'h7F90	;
				14'b00111100101010: Data_out <= 16'h7F91	;
				14'b00111100101011: Data_out <= 16'h7F92	;
				14'b00111100101100: Data_out <= 16'h7F93	;
				14'b00111100101101: Data_out <= 16'h7F94	;
				14'b00111100101110: Data_out <= 16'h7F95	;
				14'b00111100101111: Data_out <= 16'h7F96	;
				14'b00111100110000: Data_out <= 16'h7F97	;
				14'b00111100110001: Data_out <= 16'h7F98	;
				14'b00111100110010: Data_out <= 16'h7F99	;
				14'b00111100110011: Data_out <= 16'h7F9A	;
				14'b00111100110100: Data_out <= 16'h7F9B	;
				14'b00111100110101: Data_out <= 16'h7F9C	;
				14'b00111100110110: Data_out <= 16'h7F9D	;
				14'b00111100110111: Data_out <= 16'h7F9E	;
				14'b00111100111000: Data_out <= 16'h7F9F	;
				14'b00111100111001: Data_out <= 16'h7FA0	;
				14'b00111100111010: Data_out <= 16'h7FA1	;
				14'b00111100111011: Data_out <= 16'h7FA2	;
				14'b00111100111100: Data_out <= 16'h7FA3	;
				14'b00111100111101: Data_out <= 16'h7FA4	;
				14'b00111100111110: Data_out <= 16'h7FA4	;
				14'b00111100111111: Data_out <= 16'h7FA5	;
				14'b00111101000000: Data_out <= 16'h7FA6	;
				14'b00111101000001: Data_out <= 16'h7FA7	;
				14'b00111101000010: Data_out <= 16'h7FA8	;
				14'b00111101000011: Data_out <= 16'h7FA9	;
				14'b00111101000100: Data_out <= 16'h7FAA	;
				14'b00111101000101: Data_out <= 16'h7FAB	;
				14'b00111101000110: Data_out <= 16'h7FAC	;
				14'b00111101000111: Data_out <= 16'h7FAD	;
				14'b00111101001000: Data_out <= 16'h7FAE	;
				14'b00111101001001: Data_out <= 16'h7FAE	;
				14'b00111101001010: Data_out <= 16'h7FAF	;
				14'b00111101001011: Data_out <= 16'h7FB0	;
				14'b00111101001100: Data_out <= 16'h7FB1	;
				14'b00111101001101: Data_out <= 16'h7FB2	;
				14'b00111101001110: Data_out <= 16'h7FB3	;
				14'b00111101001111: Data_out <= 16'h7FB4	;
				14'b00111101010000: Data_out <= 16'h7FB4	;
				14'b00111101010001: Data_out <= 16'h7FB5	;
				14'b00111101010010: Data_out <= 16'h7FB6	;
				14'b00111101010011: Data_out <= 16'h7FB7	;
				14'b00111101010100: Data_out <= 16'h7FB8	;
				14'b00111101010101: Data_out <= 16'h7FB9	;
				14'b00111101010110: Data_out <= 16'h7FB9	;
				14'b00111101010111: Data_out <= 16'h7FBA	;
				14'b00111101011000: Data_out <= 16'h7FBB	;
				14'b00111101011001: Data_out <= 16'h7FBC	;
				14'b00111101011010: Data_out <= 16'h7FBD	;
				14'b00111101011011: Data_out <= 16'h7FBE	;
				14'b00111101011100: Data_out <= 16'h7FBE	;
				14'b00111101011101: Data_out <= 16'h7FBF	;
				14'b00111101011110: Data_out <= 16'h7FC0	;
				14'b00111101011111: Data_out <= 16'h7FC1	;
				14'b00111101100000: Data_out <= 16'h7FC1	;
				14'b00111101100001: Data_out <= 16'h7FC2	;
				14'b00111101100010: Data_out <= 16'h7FC3	;
				14'b00111101100011: Data_out <= 16'h7FC4	;
				14'b00111101100100: Data_out <= 16'h7FC4	;
				14'b00111101100101: Data_out <= 16'h7FC5	;
				14'b00111101100110: Data_out <= 16'h7FC6	;
				14'b00111101100111: Data_out <= 16'h7FC7	;
				14'b00111101101000: Data_out <= 16'h7FC7	;
				14'b00111101101001: Data_out <= 16'h7FC8	;
				14'b00111101101010: Data_out <= 16'h7FC9	;
				14'b00111101101011: Data_out <= 16'h7FCA	;
				14'b00111101101100: Data_out <= 16'h7FCA	;
				14'b00111101101101: Data_out <= 16'h7FCB	;
				14'b00111101101110: Data_out <= 16'h7FCC	;
				14'b00111101101111: Data_out <= 16'h7FCC	;
				14'b00111101110000: Data_out <= 16'h7FCD	;
				14'b00111101110001: Data_out <= 16'h7FCE	;
				14'b00111101110010: Data_out <= 16'h7FCF	;
				14'b00111101110011: Data_out <= 16'h7FCF	;
				14'b00111101110100: Data_out <= 16'h7FD0	;
				14'b00111101110101: Data_out <= 16'h7FD1	;
				14'b00111101110110: Data_out <= 16'h7FD1	;
				14'b00111101110111: Data_out <= 16'h7FD2	;
				14'b00111101111000: Data_out <= 16'h7FD3	;
				14'b00111101111001: Data_out <= 16'h7FD3	;
				14'b00111101111010: Data_out <= 16'h7FD4	;
				14'b00111101111011: Data_out <= 16'h7FD4	;
				14'b00111101111100: Data_out <= 16'h7FD5	;
				14'b00111101111101: Data_out <= 16'h7FD6	;
				14'b00111101111110: Data_out <= 16'h7FD6	;
				14'b00111101111111: Data_out <= 16'h7FD7	;
				14'b00111110000000: Data_out <= 16'h7FD8	;
				14'b00111110000001: Data_out <= 16'h7FD8	;
				14'b00111110000010: Data_out <= 16'h7FD9	;
				14'b00111110000011: Data_out <= 16'h7FD9	;
				14'b00111110000100: Data_out <= 16'h7FDA	;
				14'b00111110000101: Data_out <= 16'h7FDB	;
				14'b00111110000110: Data_out <= 16'h7FDB	;
				14'b00111110000111: Data_out <= 16'h7FDC	;
				14'b00111110001000: Data_out <= 16'h7FDC	;
				14'b00111110001001: Data_out <= 16'h7FDD	;
				14'b00111110001010: Data_out <= 16'h7FDE	;
				14'b00111110001011: Data_out <= 16'h7FDE	;
				14'b00111110001100: Data_out <= 16'h7FDF	;
				14'b00111110001101: Data_out <= 16'h7FDF	;
				14'b00111110001110: Data_out <= 16'h7FE0	;
				14'b00111110001111: Data_out <= 16'h7FE0	;
				14'b00111110010000: Data_out <= 16'h7FE1	;
				14'b00111110010001: Data_out <= 16'h7FE1	;
				14'b00111110010010: Data_out <= 16'h7FE2	;
				14'b00111110010011: Data_out <= 16'h7FE2	;
				14'b00111110010100: Data_out <= 16'h7FE3	;
				14'b00111110010101: Data_out <= 16'h7FE4	;
				14'b00111110010110: Data_out <= 16'h7FE4	;
				14'b00111110010111: Data_out <= 16'h7FE5	;
				14'b00111110011000: Data_out <= 16'h7FE5	;
				14'b00111110011001: Data_out <= 16'h7FE6	;
				14'b00111110011010: Data_out <= 16'h7FE6	;
				14'b00111110011011: Data_out <= 16'h7FE7	;
				14'b00111110011100: Data_out <= 16'h7FE7	;
				14'b00111110011101: Data_out <= 16'h7FE7	;
				14'b00111110011110: Data_out <= 16'h7FE8	;
				14'b00111110011111: Data_out <= 16'h7FE8	;
				14'b00111110100000: Data_out <= 16'h7FE9	;
				14'b00111110100001: Data_out <= 16'h7FE9	;
				14'b00111110100010: Data_out <= 16'h7FEA	;
				14'b00111110100011: Data_out <= 16'h7FEA	;
				14'b00111110100100: Data_out <= 16'h7FEB	;
				14'b00111110100101: Data_out <= 16'h7FEB	;
				14'b00111110100110: Data_out <= 16'h7FEC	;
				14'b00111110100111: Data_out <= 16'h7FEC	;
				14'b00111110101000: Data_out <= 16'h7FEC	;
				14'b00111110101001: Data_out <= 16'h7FED	;
				14'b00111110101010: Data_out <= 16'h7FED	;
				14'b00111110101011: Data_out <= 16'h7FEE	;
				14'b00111110101100: Data_out <= 16'h7FEE	;
				14'b00111110101101: Data_out <= 16'h7FEF	;
				14'b00111110101110: Data_out <= 16'h7FEF	;
				14'b00111110101111: Data_out <= 16'h7FEF	;
				14'b00111110110000: Data_out <= 16'h7FF0	;
				14'b00111110110001: Data_out <= 16'h7FF0	;
				14'b00111110110010: Data_out <= 16'h7FF0	;
				14'b00111110110011: Data_out <= 16'h7FF1	;
				14'b00111110110100: Data_out <= 16'h7FF1	;
				14'b00111110110101: Data_out <= 16'h7FF2	;
				14'b00111110110110: Data_out <= 16'h7FF2	;
				14'b00111110110111: Data_out <= 16'h7FF2	;
				14'b00111110111000: Data_out <= 16'h7FF3	;
				14'b00111110111001: Data_out <= 16'h7FF3	;
				14'b00111110111010: Data_out <= 16'h7FF3	;
				14'b00111110111011: Data_out <= 16'h7FF4	;
				14'b00111110111100: Data_out <= 16'h7FF4	;
				14'b00111110111101: Data_out <= 16'h7FF4	;
				14'b00111110111110: Data_out <= 16'h7FF5	;
				14'b00111110111111: Data_out <= 16'h7FF5	;
				14'b00111111000000: Data_out <= 16'h7FF5	;
				14'b00111111000001: Data_out <= 16'h7FF6	;
				14'b00111111000010: Data_out <= 16'h7FF6	;
				14'b00111111000011: Data_out <= 16'h7FF6	;
				14'b00111111000100: Data_out <= 16'h7FF6	;
				14'b00111111000101: Data_out <= 16'h7FF7	;
				14'b00111111000110: Data_out <= 16'h7FF7	;
				14'b00111111000111: Data_out <= 16'h7FF7	;
				14'b00111111001000: Data_out <= 16'h7FF8	;
				14'b00111111001001: Data_out <= 16'h7FF8	;
				14'b00111111001010: Data_out <= 16'h7FF8	;
				14'b00111111001011: Data_out <= 16'h7FF8	;
				14'b00111111001100: Data_out <= 16'h7FF9	;
				14'b00111111001101: Data_out <= 16'h7FF9	;
				14'b00111111001110: Data_out <= 16'h7FF9	;
				14'b00111111001111: Data_out <= 16'h7FF9	;
				14'b00111111010000: Data_out <= 16'h7FFA	;
				14'b00111111010001: Data_out <= 16'h7FFA	;
				14'b00111111010010: Data_out <= 16'h7FFA	;
				14'b00111111010011: Data_out <= 16'h7FFA	;
				14'b00111111010100: Data_out <= 16'h7FFA	;
				14'b00111111010101: Data_out <= 16'h7FFB	;
				14'b00111111010110: Data_out <= 16'h7FFB	;
				14'b00111111010111: Data_out <= 16'h7FFB	;
				14'b00111111011000: Data_out <= 16'h7FFB	;
				14'b00111111011001: Data_out <= 16'h7FFB	;
				14'b00111111011010: Data_out <= 16'h7FFC	;
				14'b00111111011011: Data_out <= 16'h7FFC	;
				14'b00111111011100: Data_out <= 16'h7FFC	;
				14'b00111111011101: Data_out <= 16'h7FFC	;
				14'b00111111011110: Data_out <= 16'h7FFC	;
				14'b00111111011111: Data_out <= 16'h7FFC	;
				14'b00111111100000: Data_out <= 16'h7FFD	;
				14'b00111111100001: Data_out <= 16'h7FFD	;
				14'b00111111100010: Data_out <= 16'h7FFD	;
				14'b00111111100011: Data_out <= 16'h7FFD	;
				14'b00111111100100: Data_out <= 16'h7FFD	;
				14'b00111111100101: Data_out <= 16'h7FFD	;
				14'b00111111100110: Data_out <= 16'h7FFD	;
				14'b00111111100111: Data_out <= 16'h7FFE	;
				14'b00111111101000: Data_out <= 16'h7FFE	;
				14'b00111111101001: Data_out <= 16'h7FFE	;
				14'b00111111101010: Data_out <= 16'h7FFE	;
				14'b00111111101011: Data_out <= 16'h7FFE	;
				14'b00111111101100: Data_out <= 16'h7FFE	;
				14'b00111111101101: Data_out <= 16'h7FFE	;
				14'b00111111101110: Data_out <= 16'h7FFE	;
				14'b00111111101111: Data_out <= 16'h7FFE	;
				14'b00111111110000: Data_out <= 16'h7FFE	;
				14'b00111111110001: Data_out <= 16'h7FFF	;
				14'b00111111110010: Data_out <= 16'h7FFF	;
				14'b00111111110011: Data_out <= 16'h7FFF	;
				14'b00111111110100: Data_out <= 16'h7FFF	;
				14'b00111111110101: Data_out <= 16'h7FFF	;
				14'b00111111110110: Data_out <= 16'h7FFF	;
				14'b00111111110111: Data_out <= 16'h7FFF	;
				14'b00111111111000: Data_out <= 16'h7FFF	;
				14'b00111111111001: Data_out <= 16'h7FFF	;
				14'b00111111111010: Data_out <= 16'h7FFF	;
				14'b00111111111011: Data_out <= 16'h7FFF	;
				14'b00111111111100: Data_out <= 16'h7FFF	;
				14'b00111111111101: Data_out <= 16'h7FFF	;
				14'b00111111111110: Data_out <= 16'h7FFF	;
				14'b00111111111111: Data_out <= 16'h7FFF	;
				/////////////////////////////////////////////////////////////////////////////////////////////
				//	posedge	half-cycle of fall......
				14'b01000000000000: Data_out <= 16'h7FFF	;
				14'b01000000000001: Data_out <= 16'h7FFF	;
				14'b01000000000010: Data_out <= 16'h7FFF	;
				14'b01000000000011: Data_out <= 16'h7FFF	;
				14'b01000000000100: Data_out <= 16'h7FFF	;
				14'b01000000000101: Data_out <= 16'h7FFF	;
				14'b01000000000110: Data_out <= 16'h7FFF	;
				14'b01000000000111: Data_out <= 16'h7FFF	;
				14'b01000000001000: Data_out <= 16'h7FFF	;
				14'b01000000001001: Data_out <= 16'h7FFF	;
				14'b01000000001010: Data_out <= 16'h7FFF	;
				14'b01000000001011: Data_out <= 16'h7FFF	;
				14'b01000000001100: Data_out <= 16'h7FFF	;
				14'b01000000001101: Data_out <= 16'h7FFF	;
				14'b01000000001110: Data_out <= 16'h7FFF	;
				14'b01000000001111: Data_out <= 16'h7FFF	;
				14'b01000000010000: Data_out <= 16'h7FFE	;
				14'b01000000010001: Data_out <= 16'h7FFE	;
				14'b01000000010010: Data_out <= 16'h7FFE	;
				14'b01000000010011: Data_out <= 16'h7FFE	;
				14'b01000000010100: Data_out <= 16'h7FFE	;
				14'b01000000010101: Data_out <= 16'h7FFE	;
				14'b01000000010110: Data_out <= 16'h7FFE	;
				14'b01000000010111: Data_out <= 16'h7FFE	;
				14'b01000000011000: Data_out <= 16'h7FFE	;
				14'b01000000011001: Data_out <= 16'h7FFE	;
				14'b01000000011010: Data_out <= 16'h7FFD	;
				14'b01000000011011: Data_out <= 16'h7FFD	;
				14'b01000000011100: Data_out <= 16'h7FFD	;
				14'b01000000011101: Data_out <= 16'h7FFD	;
				14'b01000000011110: Data_out <= 16'h7FFD	;
				14'b01000000011111: Data_out <= 16'h7FFD	;
				14'b01000000100000: Data_out <= 16'h7FFD	;
				14'b01000000100001: Data_out <= 16'h7FFC	;
				14'b01000000100010: Data_out <= 16'h7FFC	;
				14'b01000000100011: Data_out <= 16'h7FFC	;
				14'b01000000100100: Data_out <= 16'h7FFC	;
				14'b01000000100101: Data_out <= 16'h7FFC	;
				14'b01000000100110: Data_out <= 16'h7FFC	;
				14'b01000000100111: Data_out <= 16'h7FFB	;
				14'b01000000101000: Data_out <= 16'h7FFB	;
				14'b01000000101001: Data_out <= 16'h7FFB	;
				14'b01000000101010: Data_out <= 16'h7FFB	;
				14'b01000000101011: Data_out <= 16'h7FFB	;
				14'b01000000101100: Data_out <= 16'h7FFA	;
				14'b01000000101101: Data_out <= 16'h7FFA	;
				14'b01000000101110: Data_out <= 16'h7FFA	;
				14'b01000000101111: Data_out <= 16'h7FFA	;
				14'b01000000110000: Data_out <= 16'h7FFA	;
				14'b01000000110001: Data_out <= 16'h7FF9	;
				14'b01000000110010: Data_out <= 16'h7FF9	;
				14'b01000000110011: Data_out <= 16'h7FF9	;
				14'b01000000110100: Data_out <= 16'h7FF9	;
				14'b01000000110101: Data_out <= 16'h7FF8	;
				14'b01000000110110: Data_out <= 16'h7FF8	;
				14'b01000000110111: Data_out <= 16'h7FF8	;
				14'b01000000111000: Data_out <= 16'h7FF8	;
				14'b01000000111001: Data_out <= 16'h7FF7	;
				14'b01000000111010: Data_out <= 16'h7FF7	;
				14'b01000000111011: Data_out <= 16'h7FF7	;
				14'b01000000111100: Data_out <= 16'h7FF6	;
				14'b01000000111101: Data_out <= 16'h7FF6	;
				14'b01000000111110: Data_out <= 16'h7FF6	;
				14'b01000000111111: Data_out <= 16'h7FF6	;
				14'b01000001000000: Data_out <= 16'h7FF5	;
				14'b01000001000001: Data_out <= 16'h7FF5	;
				14'b01000001000010: Data_out <= 16'h7FF5	;
				14'b01000001000011: Data_out <= 16'h7FF4	;
				14'b01000001000100: Data_out <= 16'h7FF4	;
				14'b01000001000101: Data_out <= 16'h7FF4	;
				14'b01000001000110: Data_out <= 16'h7FF3	;
				14'b01000001000111: Data_out <= 16'h7FF3	;
				14'b01000001001000: Data_out <= 16'h7FF3	;
				14'b01000001001001: Data_out <= 16'h7FF2	;
				14'b01000001001010: Data_out <= 16'h7FF2	;
				14'b01000001001011: Data_out <= 16'h7FF2	;
				14'b01000001001100: Data_out <= 16'h7FF1	;
				14'b01000001001101: Data_out <= 16'h7FF1	;
				14'b01000001001110: Data_out <= 16'h7FF0	;
				14'b01000001001111: Data_out <= 16'h7FF0	;
				14'b01000001010000: Data_out <= 16'h7FF0	;
				14'b01000001010001: Data_out <= 16'h7FEF	;
				14'b01000001010010: Data_out <= 16'h7FEF	;
				14'b01000001010011: Data_out <= 16'h7FEF	;
				14'b01000001010100: Data_out <= 16'h7FEE	;
				14'b01000001010101: Data_out <= 16'h7FEE	;
				14'b01000001010110: Data_out <= 16'h7FED	;
				14'b01000001010111: Data_out <= 16'h7FED	;
				14'b01000001011000: Data_out <= 16'h7FEC	;
				14'b01000001011001: Data_out <= 16'h7FEC	;
				14'b01000001011010: Data_out <= 16'h7FEC	;
				14'b01000001011011: Data_out <= 16'h7FEB	;
				14'b01000001011100: Data_out <= 16'h7FEB	;
				14'b01000001011101: Data_out <= 16'h7FEA	;
				14'b01000001011110: Data_out <= 16'h7FEA	;
				14'b01000001011111: Data_out <= 16'h7FE9	;
				14'b01000001100000: Data_out <= 16'h7FE9	;
				14'b01000001100001: Data_out <= 16'h7FE8	;
				14'b01000001100010: Data_out <= 16'h7FE8	;
				14'b01000001100011: Data_out <= 16'h7FE7	;
				14'b01000001100100: Data_out <= 16'h7FE7	;
				14'b01000001100101: Data_out <= 16'h7FE7	;
				14'b01000001100110: Data_out <= 16'h7FE6	;
				14'b01000001100111: Data_out <= 16'h7FE6	;
				14'b01000001101000: Data_out <= 16'h7FE5	;
				14'b01000001101001: Data_out <= 16'h7FE5	;
				14'b01000001101010: Data_out <= 16'h7FE4	;
				14'b01000001101011: Data_out <= 16'h7FE4	;
				14'b01000001101100: Data_out <= 16'h7FE3	;
				14'b01000001101101: Data_out <= 16'h7FE2	;
				14'b01000001101110: Data_out <= 16'h7FE2	;
				14'b01000001101111: Data_out <= 16'h7FE1	;
				14'b01000001110000: Data_out <= 16'h7FE1	;
				14'b01000001110001: Data_out <= 16'h7FE0	;
				14'b01000001110010: Data_out <= 16'h7FE0	;
				14'b01000001110011: Data_out <= 16'h7FDF	;
				14'b01000001110100: Data_out <= 16'h7FDF	;
				14'b01000001110101: Data_out <= 16'h7FDE	;
				14'b01000001110110: Data_out <= 16'h7FDE	;
				14'b01000001110111: Data_out <= 16'h7FDD	;
				14'b01000001111000: Data_out <= 16'h7FDC	;
				14'b01000001111001: Data_out <= 16'h7FDC	;
				14'b01000001111010: Data_out <= 16'h7FDB	;
				14'b01000001111011: Data_out <= 16'h7FDB	;
				14'b01000001111100: Data_out <= 16'h7FDA	;
				14'b01000001111101: Data_out <= 16'h7FD9	;
				14'b01000001111110: Data_out <= 16'h7FD9	;
				14'b01000001111111: Data_out <= 16'h7FD8	;
				14'b01000010000000: Data_out <= 16'h7FD8	;
				14'b01000010000001: Data_out <= 16'h7FD7	;
				14'b01000010000010: Data_out <= 16'h7FD6	;
				14'b01000010000011: Data_out <= 16'h7FD6	;
				14'b01000010000100: Data_out <= 16'h7FD5	;
				14'b01000010000101: Data_out <= 16'h7FD4	;
				14'b01000010000110: Data_out <= 16'h7FD4	;
				14'b01000010000111: Data_out <= 16'h7FD3	;
				14'b01000010001000: Data_out <= 16'h7FD3	;
				14'b01000010001001: Data_out <= 16'h7FD2	;
				14'b01000010001010: Data_out <= 16'h7FD1	;
				14'b01000010001011: Data_out <= 16'h7FD1	;
				14'b01000010001100: Data_out <= 16'h7FD0	;
				14'b01000010001101: Data_out <= 16'h7FCF	;
				14'b01000010001110: Data_out <= 16'h7FCF	;
				14'b01000010001111: Data_out <= 16'h7FCE	;
				14'b01000010010000: Data_out <= 16'h7FCD	;
				14'b01000010010001: Data_out <= 16'h7FCC	;
				14'b01000010010010: Data_out <= 16'h7FCC	;
				14'b01000010010011: Data_out <= 16'h7FCB	;
				14'b01000010010100: Data_out <= 16'h7FCA	;
				14'b01000010010101: Data_out <= 16'h7FCA	;
				14'b01000010010110: Data_out <= 16'h7FC9	;
				14'b01000010010111: Data_out <= 16'h7FC8	;
				14'b01000010011000: Data_out <= 16'h7FC7	;
				14'b01000010011001: Data_out <= 16'h7FC7	;
				14'b01000010011010: Data_out <= 16'h7FC6	;
				14'b01000010011011: Data_out <= 16'h7FC5	;
				14'b01000010011100: Data_out <= 16'h7FC4	;
				14'b01000010011101: Data_out <= 16'h7FC4	;
				14'b01000010011110: Data_out <= 16'h7FC3	;
				14'b01000010011111: Data_out <= 16'h7FC2	;
				14'b01000010100000: Data_out <= 16'h7FC1	;
				14'b01000010100001: Data_out <= 16'h7FC1	;
				14'b01000010100010: Data_out <= 16'h7FC0	;
				14'b01000010100011: Data_out <= 16'h7FBF	;
				14'b01000010100100: Data_out <= 16'h7FBE	;
				14'b01000010100101: Data_out <= 16'h7FBE	;
				14'b01000010100110: Data_out <= 16'h7FBD	;
				14'b01000010100111: Data_out <= 16'h7FBC	;
				14'b01000010101000: Data_out <= 16'h7FBB	;
				14'b01000010101001: Data_out <= 16'h7FBA	;
				14'b01000010101010: Data_out <= 16'h7FB9	;
				14'b01000010101011: Data_out <= 16'h7FB9	;
				14'b01000010101100: Data_out <= 16'h7FB8	;
				14'b01000010101101: Data_out <= 16'h7FB7	;
				14'b01000010101110: Data_out <= 16'h7FB6	;
				14'b01000010101111: Data_out <= 16'h7FB5	;
				14'b01000010110000: Data_out <= 16'h7FB4	;
				14'b01000010110001: Data_out <= 16'h7FB4	;
				14'b01000010110010: Data_out <= 16'h7FB3	;
				14'b01000010110011: Data_out <= 16'h7FB2	;
				14'b01000010110100: Data_out <= 16'h7FB1	;
				14'b01000010110101: Data_out <= 16'h7FB0	;
				14'b01000010110110: Data_out <= 16'h7FAF	;
				14'b01000010110111: Data_out <= 16'h7FAE	;
				14'b01000010111000: Data_out <= 16'h7FAE	;
				14'b01000010111001: Data_out <= 16'h7FAD	;
				14'b01000010111010: Data_out <= 16'h7FAC	;
				14'b01000010111011: Data_out <= 16'h7FAB	;
				14'b01000010111100: Data_out <= 16'h7FAA	;
				14'b01000010111101: Data_out <= 16'h7FA9	;
				14'b01000010111110: Data_out <= 16'h7FA8	;
				14'b01000010111111: Data_out <= 16'h7FA7	;
				14'b01000011000000: Data_out <= 16'h7FA6	;
				14'b01000011000001: Data_out <= 16'h7FA5	;
				14'b01000011000010: Data_out <= 16'h7FA4	;
				14'b01000011000011: Data_out <= 16'h7FA4	;
				14'b01000011000100: Data_out <= 16'h7FA3	;
				14'b01000011000101: Data_out <= 16'h7FA2	;
				14'b01000011000110: Data_out <= 16'h7FA1	;
				14'b01000011000111: Data_out <= 16'h7FA0	;
				14'b01000011001000: Data_out <= 16'h7F9F	;
				14'b01000011001001: Data_out <= 16'h7F9E	;
				14'b01000011001010: Data_out <= 16'h7F9D	;
				14'b01000011001011: Data_out <= 16'h7F9C	;
				14'b01000011001100: Data_out <= 16'h7F9B	;
				14'b01000011001101: Data_out <= 16'h7F9A	;
				14'b01000011001110: Data_out <= 16'h7F99	;
				14'b01000011001111: Data_out <= 16'h7F98	;
				14'b01000011010000: Data_out <= 16'h7F97	;
				14'b01000011010001: Data_out <= 16'h7F96	;
				14'b01000011010010: Data_out <= 16'h7F95	;
				14'b01000011010011: Data_out <= 16'h7F94	;
				14'b01000011010100: Data_out <= 16'h7F93	;
				14'b01000011010101: Data_out <= 16'h7F92	;
				14'b01000011010110: Data_out <= 16'h7F91	;
				14'b01000011010111: Data_out <= 16'h7F90	;
				14'b01000011011000: Data_out <= 16'h7F8F	;
				14'b01000011011001: Data_out <= 16'h7F8E	;
				14'b01000011011010: Data_out <= 16'h7F8D	;
				14'b01000011011011: Data_out <= 16'h7F8C	;
				14'b01000011011100: Data_out <= 16'h7F8B	;
				14'b01000011011101: Data_out <= 16'h7F89	;
				14'b01000011011110: Data_out <= 16'h7F88	;
				14'b01000011011111: Data_out <= 16'h7F87	;
				14'b01000011100000: Data_out <= 16'h7F86	;
				14'b01000011100001: Data_out <= 16'h7F85	;
				14'b01000011100010: Data_out <= 16'h7F84	;
				14'b01000011100011: Data_out <= 16'h7F83	;
				14'b01000011100100: Data_out <= 16'h7F82	;
				14'b01000011100101: Data_out <= 16'h7F81	;
				14'b01000011100110: Data_out <= 16'h7F80	;
				14'b01000011100111: Data_out <= 16'h7F7F	;
				14'b01000011101000: Data_out <= 16'h7F7D	;
				14'b01000011101001: Data_out <= 16'h7F7C	;
				14'b01000011101010: Data_out <= 16'h7F7B	;
				14'b01000011101011: Data_out <= 16'h7F7A	;
				14'b01000011101100: Data_out <= 16'h7F79	;
				14'b01000011101101: Data_out <= 16'h7F78	;
				14'b01000011101110: Data_out <= 16'h7F77	;
				14'b01000011101111: Data_out <= 16'h7F76	;
				14'b01000011110000: Data_out <= 16'h7F74	;
				14'b01000011110001: Data_out <= 16'h7F73	;
				14'b01000011110010: Data_out <= 16'h7F72	;
				14'b01000011110011: Data_out <= 16'h7F71	;
				14'b01000011110100: Data_out <= 16'h7F70	;
				14'b01000011110101: Data_out <= 16'h7F6F	;
				14'b01000011110110: Data_out <= 16'h7F6D	;
				14'b01000011110111: Data_out <= 16'h7F6C	;
				14'b01000011111000: Data_out <= 16'h7F6B	;
				14'b01000011111001: Data_out <= 16'h7F6A	;
				14'b01000011111010: Data_out <= 16'h7F69	;
				14'b01000011111011: Data_out <= 16'h7F67	;
				14'b01000011111100: Data_out <= 16'h7F66	;
				14'b01000011111101: Data_out <= 16'h7F65	;
				14'b01000011111110: Data_out <= 16'h7F64	;
				14'b01000011111111: Data_out <= 16'h7F63	;
				14'b01000100000000: Data_out <= 16'h7F61	;
				14'b01000100000001: Data_out <= 16'h7F60	;
				14'b01000100000010: Data_out <= 16'h7F5F	;
				14'b01000100000011: Data_out <= 16'h7F5E	;
				14'b01000100000100: Data_out <= 16'h7F5C	;
				14'b01000100000101: Data_out <= 16'h7F5B	;
				14'b01000100000110: Data_out <= 16'h7F5A	;
				14'b01000100000111: Data_out <= 16'h7F59	;
				14'b01000100001000: Data_out <= 16'h7F57	;
				14'b01000100001001: Data_out <= 16'h7F56	;
				14'b01000100001010: Data_out <= 16'h7F55	;
				14'b01000100001011: Data_out <= 16'h7F53	;
				14'b01000100001100: Data_out <= 16'h7F52	;
				14'b01000100001101: Data_out <= 16'h7F51	;
				14'b01000100001110: Data_out <= 16'h7F50	;
				14'b01000100001111: Data_out <= 16'h7F4E	;
				14'b01000100010000: Data_out <= 16'h7F4D	;
				14'b01000100010001: Data_out <= 16'h7F4C	;
				14'b01000100010010: Data_out <= 16'h7F4A	;
				14'b01000100010011: Data_out <= 16'h7F49	;
				14'b01000100010100: Data_out <= 16'h7F48	;
				14'b01000100010101: Data_out <= 16'h7F46	;
				14'b01000100010110: Data_out <= 16'h7F45	;
				14'b01000100010111: Data_out <= 16'h7F44	;
				14'b01000100011000: Data_out <= 16'h7F42	;
				14'b01000100011001: Data_out <= 16'h7F41	;
				14'b01000100011010: Data_out <= 16'h7F40	;
				14'b01000100011011: Data_out <= 16'h7F3E	;
				14'b01000100011100: Data_out <= 16'h7F3D	;
				14'b01000100011101: Data_out <= 16'h7F3C	;
				14'b01000100011110: Data_out <= 16'h7F3A	;
				14'b01000100011111: Data_out <= 16'h7F39	;
				14'b01000100100000: Data_out <= 16'h7F37	;
				14'b01000100100001: Data_out <= 16'h7F36	;
				14'b01000100100010: Data_out <= 16'h7F35	;
				14'b01000100100011: Data_out <= 16'h7F33	;
				14'b01000100100100: Data_out <= 16'h7F32	;
				14'b01000100100101: Data_out <= 16'h7F30	;
				14'b01000100100110: Data_out <= 16'h7F2F	;
				14'b01000100100111: Data_out <= 16'h7F2E	;
				14'b01000100101000: Data_out <= 16'h7F2C	;
				14'b01000100101001: Data_out <= 16'h7F2B	;
				14'b01000100101010: Data_out <= 16'h7F29	;
				14'b01000100101011: Data_out <= 16'h7F28	;
				14'b01000100101100: Data_out <= 16'h7F26	;
				14'b01000100101101: Data_out <= 16'h7F25	;
				14'b01000100101110: Data_out <= 16'h7F24	;
				14'b01000100101111: Data_out <= 16'h7F22	;
				14'b01000100110000: Data_out <= 16'h7F21	;
				14'b01000100110001: Data_out <= 16'h7F1F	;
				14'b01000100110010: Data_out <= 16'h7F1E	;
				14'b01000100110011: Data_out <= 16'h7F1C	;
				14'b01000100110100: Data_out <= 16'h7F1B	;
				14'b01000100110101: Data_out <= 16'h7F19	;
				14'b01000100110110: Data_out <= 16'h7F18	;
				14'b01000100110111: Data_out <= 16'h7F16	;
				14'b01000100111000: Data_out <= 16'h7F15	;
				14'b01000100111001: Data_out <= 16'h7F13	;
				14'b01000100111010: Data_out <= 16'h7F12	;
				14'b01000100111011: Data_out <= 16'h7F10	;
				14'b01000100111100: Data_out <= 16'h7F0F	;
				14'b01000100111101: Data_out <= 16'h7F0D	;
				14'b01000100111110: Data_out <= 16'h7F0C	;
				14'b01000100111111: Data_out <= 16'h7F0A	;
				14'b01000101000000: Data_out <= 16'h7F09	;
				14'b01000101000001: Data_out <= 16'h7F07	;
				14'b01000101000010: Data_out <= 16'h7F06	;
				14'b01000101000011: Data_out <= 16'h7F04	;
				14'b01000101000100: Data_out <= 16'h7F02	;
				14'b01000101000101: Data_out <= 16'h7F01	;
				14'b01000101000110: Data_out <= 16'h7EFF	;
				14'b01000101000111: Data_out <= 16'h7EFE	;
				14'b01000101001000: Data_out <= 16'h7EFC	;
				14'b01000101001001: Data_out <= 16'h7EFB	;
				14'b01000101001010: Data_out <= 16'h7EF9	;
				14'b01000101001011: Data_out <= 16'h7EF7	;
				14'b01000101001100: Data_out <= 16'h7EF6	;
				14'b01000101001101: Data_out <= 16'h7EF4	;
				14'b01000101001110: Data_out <= 16'h7EF3	;
				14'b01000101001111: Data_out <= 16'h7EF1	;
				14'b01000101010000: Data_out <= 16'h7EEF	;
				14'b01000101010001: Data_out <= 16'h7EEE	;
				14'b01000101010010: Data_out <= 16'h7EEC	;
				14'b01000101010011: Data_out <= 16'h7EEB	;
				14'b01000101010100: Data_out <= 16'h7EE9	;
				14'b01000101010101: Data_out <= 16'h7EE7	;
				14'b01000101010110: Data_out <= 16'h7EE6	;
				14'b01000101010111: Data_out <= 16'h7EE4	;
				14'b01000101011000: Data_out <= 16'h7EE2	;
				14'b01000101011001: Data_out <= 16'h7EE1	;
				14'b01000101011010: Data_out <= 16'h7EDF	;
				14'b01000101011011: Data_out <= 16'h7EDD	;
				14'b01000101011100: Data_out <= 16'h7EDC	;
				14'b01000101011101: Data_out <= 16'h7EDA	;
				14'b01000101011110: Data_out <= 16'h7ED8	;
				14'b01000101011111: Data_out <= 16'h7ED7	;
				14'b01000101100000: Data_out <= 16'h7ED5	;
				14'b01000101100001: Data_out <= 16'h7ED3	;
				14'b01000101100010: Data_out <= 16'h7ED2	;
				14'b01000101100011: Data_out <= 16'h7ED0	;
				14'b01000101100100: Data_out <= 16'h7ECE	;
				14'b01000101100101: Data_out <= 16'h7ECC	;
				14'b01000101100110: Data_out <= 16'h7ECB	;
				14'b01000101100111: Data_out <= 16'h7EC9	;
				14'b01000101101000: Data_out <= 16'h7EC7	;
				14'b01000101101001: Data_out <= 16'h7EC6	;
				14'b01000101101010: Data_out <= 16'h7EC4	;
				14'b01000101101011: Data_out <= 16'h7EC2	;
				14'b01000101101100: Data_out <= 16'h7EC0	;
				14'b01000101101101: Data_out <= 16'h7EBF	;
				14'b01000101101110: Data_out <= 16'h7EBD	;
				14'b01000101101111: Data_out <= 16'h7EBB	;
				14'b01000101110000: Data_out <= 16'h7EB9	;
				14'b01000101110001: Data_out <= 16'h7EB8	;
				14'b01000101110010: Data_out <= 16'h7EB6	;
				14'b01000101110011: Data_out <= 16'h7EB4	;
				14'b01000101110100: Data_out <= 16'h7EB2	;
				14'b01000101110101: Data_out <= 16'h7EB0	;
				14'b01000101110110: Data_out <= 16'h7EAF	;
				14'b01000101110111: Data_out <= 16'h7EAD	;
				14'b01000101111000: Data_out <= 16'h7EAB	;
				14'b01000101111001: Data_out <= 16'h7EA9	;
				14'b01000101111010: Data_out <= 16'h7EA7	;
				14'b01000101111011: Data_out <= 16'h7EA6	;
				14'b01000101111100: Data_out <= 16'h7EA4	;
				14'b01000101111101: Data_out <= 16'h7EA2	;
				14'b01000101111110: Data_out <= 16'h7EA0	;
				14'b01000101111111: Data_out <= 16'h7E9E	;
				14'b01000110000000: Data_out <= 16'h7E9C	;
				14'b01000110000001: Data_out <= 16'h7E9B	;
				14'b01000110000010: Data_out <= 16'h7E99	;
				14'b01000110000011: Data_out <= 16'h7E97	;
				14'b01000110000100: Data_out <= 16'h7E95	;
				14'b01000110000101: Data_out <= 16'h7E93	;
				14'b01000110000110: Data_out <= 16'h7E91	;
				14'b01000110000111: Data_out <= 16'h7E8F	;
				14'b01000110001000: Data_out <= 16'h7E8E	;
				14'b01000110001001: Data_out <= 16'h7E8C	;
				14'b01000110001010: Data_out <= 16'h7E8A	;
				14'b01000110001011: Data_out <= 16'h7E88	;
				14'b01000110001100: Data_out <= 16'h7E86	;
				14'b01000110001101: Data_out <= 16'h7E84	;
				14'b01000110001110: Data_out <= 16'h7E82	;
				14'b01000110001111: Data_out <= 16'h7E80	;
				14'b01000110010000: Data_out <= 16'h7E7E	;
				14'b01000110010001: Data_out <= 16'h7E7C	;
				14'b01000110010010: Data_out <= 16'h7E7A	;
				14'b01000110010011: Data_out <= 16'h7E79	;
				14'b01000110010100: Data_out <= 16'h7E77	;
				14'b01000110010101: Data_out <= 16'h7E75	;
				14'b01000110010110: Data_out <= 16'h7E73	;
				14'b01000110010111: Data_out <= 16'h7E71	;
				14'b01000110011000: Data_out <= 16'h7E6F	;
				14'b01000110011001: Data_out <= 16'h7E6D	;
				14'b01000110011010: Data_out <= 16'h7E6B	;
				14'b01000110011011: Data_out <= 16'h7E69	;
				14'b01000110011100: Data_out <= 16'h7E67	;
				14'b01000110011101: Data_out <= 16'h7E65	;
				14'b01000110011110: Data_out <= 16'h7E63	;
				14'b01000110011111: Data_out <= 16'h7E61	;
				14'b01000110100000: Data_out <= 16'h7E5F	;
				14'b01000110100001: Data_out <= 16'h7E5D	;
				14'b01000110100010: Data_out <= 16'h7E5B	;
				14'b01000110100011: Data_out <= 16'h7E59	;
				14'b01000110100100: Data_out <= 16'h7E57	;
				14'b01000110100101: Data_out <= 16'h7E55	;
				14'b01000110100110: Data_out <= 16'h7E53	;
				14'b01000110100111: Data_out <= 16'h7E51	;
				14'b01000110101000: Data_out <= 16'h7E4F	;
				14'b01000110101001: Data_out <= 16'h7E4D	;
				14'b01000110101010: Data_out <= 16'h7E4B	;
				14'b01000110101011: Data_out <= 16'h7E49	;
				14'b01000110101100: Data_out <= 16'h7E47	;
				14'b01000110101101: Data_out <= 16'h7E45	;
				14'b01000110101110: Data_out <= 16'h7E43	;
				14'b01000110101111: Data_out <= 16'h7E41	;
				14'b01000110110000: Data_out <= 16'h7E3E	;
				14'b01000110110001: Data_out <= 16'h7E3C	;
				14'b01000110110010: Data_out <= 16'h7E3A	;
				14'b01000110110011: Data_out <= 16'h7E38	;
				14'b01000110110100: Data_out <= 16'h7E36	;
				14'b01000110110101: Data_out <= 16'h7E34	;
				14'b01000110110110: Data_out <= 16'h7E32	;
				14'b01000110110111: Data_out <= 16'h7E30	;
				14'b01000110111000: Data_out <= 16'h7E2E	;
				14'b01000110111001: Data_out <= 16'h7E2C	;
				14'b01000110111010: Data_out <= 16'h7E29	;
				14'b01000110111011: Data_out <= 16'h7E27	;
				14'b01000110111100: Data_out <= 16'h7E25	;
				14'b01000110111101: Data_out <= 16'h7E23	;
				14'b01000110111110: Data_out <= 16'h7E21	;
				14'b01000110111111: Data_out <= 16'h7E1F	;
				14'b01000111000000: Data_out <= 16'h7E1D	;
				14'b01000111000001: Data_out <= 16'h7E1B	;
				14'b01000111000010: Data_out <= 16'h7E18	;
				14'b01000111000011: Data_out <= 16'h7E16	;
				14'b01000111000100: Data_out <= 16'h7E14	;
				14'b01000111000101: Data_out <= 16'h7E12	;
				14'b01000111000110: Data_out <= 16'h7E10	;
				14'b01000111000111: Data_out <= 16'h7E0E	;
				14'b01000111001000: Data_out <= 16'h7E0B	;
				14'b01000111001001: Data_out <= 16'h7E09	;
				14'b01000111001010: Data_out <= 16'h7E07	;
				14'b01000111001011: Data_out <= 16'h7E05	;
				14'b01000111001100: Data_out <= 16'h7E03	;
				14'b01000111001101: Data_out <= 16'h7E00	;
				14'b01000111001110: Data_out <= 16'h7DFE	;
				14'b01000111001111: Data_out <= 16'h7DFC	;
				14'b01000111010000: Data_out <= 16'h7DFA	;
				14'b01000111010001: Data_out <= 16'h7DF7	;
				14'b01000111010010: Data_out <= 16'h7DF5	;
				14'b01000111010011: Data_out <= 16'h7DF3	;
				14'b01000111010100: Data_out <= 16'h7DF1	;
				14'b01000111010101: Data_out <= 16'h7DEF	;
				14'b01000111010110: Data_out <= 16'h7DEC	;
				14'b01000111010111: Data_out <= 16'h7DEA	;
				14'b01000111011000: Data_out <= 16'h7DE8	;
				14'b01000111011001: Data_out <= 16'h7DE6	;
				14'b01000111011010: Data_out <= 16'h7DE3	;
				14'b01000111011011: Data_out <= 16'h7DE1	;
				14'b01000111011100: Data_out <= 16'h7DDF	;
				14'b01000111011101: Data_out <= 16'h7DDC	;
				14'b01000111011110: Data_out <= 16'h7DDA	;
				14'b01000111011111: Data_out <= 16'h7DD8	;
				14'b01000111100000: Data_out <= 16'h7DD6	;
				14'b01000111100001: Data_out <= 16'h7DD3	;
				14'b01000111100010: Data_out <= 16'h7DD1	;
				14'b01000111100011: Data_out <= 16'h7DCF	;
				14'b01000111100100: Data_out <= 16'h7DCC	;
				14'b01000111100101: Data_out <= 16'h7DCA	;
				14'b01000111100110: Data_out <= 16'h7DC8	;
				14'b01000111100111: Data_out <= 16'h7DC5	;
				14'b01000111101000: Data_out <= 16'h7DC3	;
				14'b01000111101001: Data_out <= 16'h7DC1	;
				14'b01000111101010: Data_out <= 16'h7DBE	;
				14'b01000111101011: Data_out <= 16'h7DBC	;
				14'b01000111101100: Data_out <= 16'h7DBA	;
				14'b01000111101101: Data_out <= 16'h7DB7	;
				14'b01000111101110: Data_out <= 16'h7DB5	;
				14'b01000111101111: Data_out <= 16'h7DB2	;
				14'b01000111110000: Data_out <= 16'h7DB0	;
				14'b01000111110001: Data_out <= 16'h7DAE	;
				14'b01000111110010: Data_out <= 16'h7DAB	;
				14'b01000111110011: Data_out <= 16'h7DA9	;
				14'b01000111110100: Data_out <= 16'h7DA7	;
				14'b01000111110101: Data_out <= 16'h7DA4	;
				14'b01000111110110: Data_out <= 16'h7DA2	;
				14'b01000111110111: Data_out <= 16'h7D9F	;
				14'b01000111111000: Data_out <= 16'h7D9D	;
				14'b01000111111001: Data_out <= 16'h7D9B	;
				14'b01000111111010: Data_out <= 16'h7D98	;
				14'b01000111111011: Data_out <= 16'h7D96	;
				14'b01000111111100: Data_out <= 16'h7D93	;
				14'b01000111111101: Data_out <= 16'h7D91	;
				14'b01000111111110: Data_out <= 16'h7D8E	;
				14'b01000111111111: Data_out <= 16'h7D8C	;
				14'b01001000000000: Data_out <= 16'h7D89	;
				14'b01001000000001: Data_out <= 16'h7D87	;
				14'b01001000000010: Data_out <= 16'h7D85	;
				14'b01001000000011: Data_out <= 16'h7D82	;
				14'b01001000000100: Data_out <= 16'h7D80	;
				14'b01001000000101: Data_out <= 16'h7D7D	;
				14'b01001000000110: Data_out <= 16'h7D7B	;
				14'b01001000000111: Data_out <= 16'h7D78	;
				14'b01001000001000: Data_out <= 16'h7D76	;
				14'b01001000001001: Data_out <= 16'h7D73	;
				14'b01001000001010: Data_out <= 16'h7D71	;
				14'b01001000001011: Data_out <= 16'h7D6E	;
				14'b01001000001100: Data_out <= 16'h7D6C	;
				14'b01001000001101: Data_out <= 16'h7D69	;
				14'b01001000001110: Data_out <= 16'h7D67	;
				14'b01001000001111: Data_out <= 16'h7D64	;
				14'b01001000010000: Data_out <= 16'h7D62	;
				14'b01001000010001: Data_out <= 16'h7D5F	;
				14'b01001000010010: Data_out <= 16'h7D5D	;
				14'b01001000010011: Data_out <= 16'h7D5A	;
				14'b01001000010100: Data_out <= 16'h7D58	;
				14'b01001000010101: Data_out <= 16'h7D55	;
				14'b01001000010110: Data_out <= 16'h7D52	;
				14'b01001000010111: Data_out <= 16'h7D50	;
				14'b01001000011000: Data_out <= 16'h7D4D	;
				14'b01001000011001: Data_out <= 16'h7D4B	;
				14'b01001000011010: Data_out <= 16'h7D48	;
				14'b01001000011011: Data_out <= 16'h7D46	;
				14'b01001000011100: Data_out <= 16'h7D43	;
				14'b01001000011101: Data_out <= 16'h7D40	;
				14'b01001000011110: Data_out <= 16'h7D3E	;
				14'b01001000011111: Data_out <= 16'h7D3B	;
				14'b01001000100000: Data_out <= 16'h7D39	;
				14'b01001000100001: Data_out <= 16'h7D36	;
				14'b01001000100010: Data_out <= 16'h7D33	;
				14'b01001000100011: Data_out <= 16'h7D31	;
				14'b01001000100100: Data_out <= 16'h7D2E	;
				14'b01001000100101: Data_out <= 16'h7D2C	;
				14'b01001000100110: Data_out <= 16'h7D29	;
				14'b01001000100111: Data_out <= 16'h7D26	;
				14'b01001000101000: Data_out <= 16'h7D24	;
				14'b01001000101001: Data_out <= 16'h7D21	;
				14'b01001000101010: Data_out <= 16'h7D1E	;
				14'b01001000101011: Data_out <= 16'h7D1C	;
				14'b01001000101100: Data_out <= 16'h7D19	;
				14'b01001000101101: Data_out <= 16'h7D16	;
				14'b01001000101110: Data_out <= 16'h7D14	;
				14'b01001000101111: Data_out <= 16'h7D11	;
				14'b01001000110000: Data_out <= 16'h7D0E	;
				14'b01001000110001: Data_out <= 16'h7D0C	;
				14'b01001000110010: Data_out <= 16'h7D09	;
				14'b01001000110011: Data_out <= 16'h7D06	;
				14'b01001000110100: Data_out <= 16'h7D04	;
				14'b01001000110101: Data_out <= 16'h7D01	;
				14'b01001000110110: Data_out <= 16'h7CFE	;
				14'b01001000110111: Data_out <= 16'h7CFC	;
				14'b01001000111000: Data_out <= 16'h7CF9	;
				14'b01001000111001: Data_out <= 16'h7CF6	;
				14'b01001000111010: Data_out <= 16'h7CF3	;
				14'b01001000111011: Data_out <= 16'h7CF1	;
				14'b01001000111100: Data_out <= 16'h7CEE	;
				14'b01001000111101: Data_out <= 16'h7CEB	;
				14'b01001000111110: Data_out <= 16'h7CE8	;
				14'b01001000111111: Data_out <= 16'h7CE6	;
				14'b01001001000000: Data_out <= 16'h7CE3	;
				14'b01001001000001: Data_out <= 16'h7CE0	;
				14'b01001001000010: Data_out <= 16'h7CDD	;
				14'b01001001000011: Data_out <= 16'h7CDB	;
				14'b01001001000100: Data_out <= 16'h7CD8	;
				14'b01001001000101: Data_out <= 16'h7CD5	;
				14'b01001001000110: Data_out <= 16'h7CD2	;
				14'b01001001000111: Data_out <= 16'h7CD0	;
				14'b01001001001000: Data_out <= 16'h7CCD	;
				14'b01001001001001: Data_out <= 16'h7CCA	;
				14'b01001001001010: Data_out <= 16'h7CC7	;
				14'b01001001001011: Data_out <= 16'h7CC4	;
				14'b01001001001100: Data_out <= 16'h7CC2	;
				14'b01001001001101: Data_out <= 16'h7CBF	;
				14'b01001001001110: Data_out <= 16'h7CBC	;
				14'b01001001001111: Data_out <= 16'h7CB9	;
				14'b01001001010000: Data_out <= 16'h7CB6	;
				14'b01001001010001: Data_out <= 16'h7CB3	;
				14'b01001001010010: Data_out <= 16'h7CB1	;
				14'b01001001010011: Data_out <= 16'h7CAE	;
				14'b01001001010100: Data_out <= 16'h7CAB	;
				14'b01001001010101: Data_out <= 16'h7CA8	;
				14'b01001001010110: Data_out <= 16'h7CA5	;
				14'b01001001010111: Data_out <= 16'h7CA2	;
				14'b01001001011000: Data_out <= 16'h7CA0	;
				14'b01001001011001: Data_out <= 16'h7C9D	;
				14'b01001001011010: Data_out <= 16'h7C9A	;
				14'b01001001011011: Data_out <= 16'h7C97	;
				14'b01001001011100: Data_out <= 16'h7C94	;
				14'b01001001011101: Data_out <= 16'h7C91	;
				14'b01001001011110: Data_out <= 16'h7C8E	;
				14'b01001001011111: Data_out <= 16'h7C8B	;
				14'b01001001100000: Data_out <= 16'h7C88	;
				14'b01001001100001: Data_out <= 16'h7C86	;
				14'b01001001100010: Data_out <= 16'h7C83	;
				14'b01001001100011: Data_out <= 16'h7C80	;
				14'b01001001100100: Data_out <= 16'h7C7D	;
				14'b01001001100101: Data_out <= 16'h7C7A	;
				14'b01001001100110: Data_out <= 16'h7C77	;
				14'b01001001100111: Data_out <= 16'h7C74	;
				14'b01001001101000: Data_out <= 16'h7C71	;
				14'b01001001101001: Data_out <= 16'h7C6E	;
				14'b01001001101010: Data_out <= 16'h7C6B	;
				14'b01001001101011: Data_out <= 16'h7C68	;
				14'b01001001101100: Data_out <= 16'h7C65	;
				14'b01001001101101: Data_out <= 16'h7C62	;
				14'b01001001101110: Data_out <= 16'h7C5F	;
				14'b01001001101111: Data_out <= 16'h7C5C	;
				14'b01001001110000: Data_out <= 16'h7C59	;
				14'b01001001110001: Data_out <= 16'h7C56	;
				14'b01001001110010: Data_out <= 16'h7C53	;
				14'b01001001110011: Data_out <= 16'h7C50	;
				14'b01001001110100: Data_out <= 16'h7C4D	;
				14'b01001001110101: Data_out <= 16'h7C4A	;
				14'b01001001110110: Data_out <= 16'h7C47	;
				14'b01001001110111: Data_out <= 16'h7C44	;
				14'b01001001111000: Data_out <= 16'h7C41	;
				14'b01001001111001: Data_out <= 16'h7C3E	;
				14'b01001001111010: Data_out <= 16'h7C3B	;
				14'b01001001111011: Data_out <= 16'h7C38	;
				14'b01001001111100: Data_out <= 16'h7C35	;
				14'b01001001111101: Data_out <= 16'h7C32	;
				14'b01001001111110: Data_out <= 16'h7C2F	;
				14'b01001001111111: Data_out <= 16'h7C2C	;
				14'b01001010000000: Data_out <= 16'h7C29	;
				14'b01001010000001: Data_out <= 16'h7C26	;
				14'b01001010000010: Data_out <= 16'h7C23	;
				14'b01001010000011: Data_out <= 16'h7C20	;
				14'b01001010000100: Data_out <= 16'h7C1D	;
				14'b01001010000101: Data_out <= 16'h7C1A	;
				14'b01001010000110: Data_out <= 16'h7C17	;
				14'b01001010000111: Data_out <= 16'h7C14	;
				14'b01001010001000: Data_out <= 16'h7C11	;
				14'b01001010001001: Data_out <= 16'h7C0D	;
				14'b01001010001010: Data_out <= 16'h7C0A	;
				14'b01001010001011: Data_out <= 16'h7C07	;
				14'b01001010001100: Data_out <= 16'h7C04	;
				14'b01001010001101: Data_out <= 16'h7C01	;
				14'b01001010001110: Data_out <= 16'h7BFE	;
				14'b01001010001111: Data_out <= 16'h7BFB	;
				14'b01001010010000: Data_out <= 16'h7BF8	;
				14'b01001010010001: Data_out <= 16'h7BF5	;
				14'b01001010010010: Data_out <= 16'h7BF1	;
				14'b01001010010011: Data_out <= 16'h7BEE	;
				14'b01001010010100: Data_out <= 16'h7BEB	;
				14'b01001010010101: Data_out <= 16'h7BE8	;
				14'b01001010010110: Data_out <= 16'h7BE5	;
				14'b01001010010111: Data_out <= 16'h7BE2	;
				14'b01001010011000: Data_out <= 16'h7BDE	;
				14'b01001010011001: Data_out <= 16'h7BDB	;
				14'b01001010011010: Data_out <= 16'h7BD8	;
				14'b01001010011011: Data_out <= 16'h7BD5	;
				14'b01001010011100: Data_out <= 16'h7BD2	;
				14'b01001010011101: Data_out <= 16'h7BCF	;
				14'b01001010011110: Data_out <= 16'h7BCB	;
				14'b01001010011111: Data_out <= 16'h7BC8	;
				14'b01001010100000: Data_out <= 16'h7BC5	;
				14'b01001010100001: Data_out <= 16'h7BC2	;
				14'b01001010100010: Data_out <= 16'h7BBF	;
				14'b01001010100011: Data_out <= 16'h7BBB	;
				14'b01001010100100: Data_out <= 16'h7BB8	;
				14'b01001010100101: Data_out <= 16'h7BB5	;
				14'b01001010100110: Data_out <= 16'h7BB2	;
				14'b01001010100111: Data_out <= 16'h7BAE	;
				14'b01001010101000: Data_out <= 16'h7BAB	;
				14'b01001010101001: Data_out <= 16'h7BA8	;
				14'b01001010101010: Data_out <= 16'h7BA5	;
				14'b01001010101011: Data_out <= 16'h7BA2	;
				14'b01001010101100: Data_out <= 16'h7B9E	;
				14'b01001010101101: Data_out <= 16'h7B9B	;
				14'b01001010101110: Data_out <= 16'h7B98	;
				14'b01001010101111: Data_out <= 16'h7B94	;
				14'b01001010110000: Data_out <= 16'h7B91	;
				14'b01001010110001: Data_out <= 16'h7B8E	;
				14'b01001010110010: Data_out <= 16'h7B8B	;
				14'b01001010110011: Data_out <= 16'h7B87	;
				14'b01001010110100: Data_out <= 16'h7B84	;
				14'b01001010110101: Data_out <= 16'h7B81	;
				14'b01001010110110: Data_out <= 16'h7B7D	;
				14'b01001010110111: Data_out <= 16'h7B7A	;
				14'b01001010111000: Data_out <= 16'h7B77	;
				14'b01001010111001: Data_out <= 16'h7B73	;
				14'b01001010111010: Data_out <= 16'h7B70	;
				14'b01001010111011: Data_out <= 16'h7B6D	;
				14'b01001010111100: Data_out <= 16'h7B6A	;
				14'b01001010111101: Data_out <= 16'h7B66	;
				14'b01001010111110: Data_out <= 16'h7B63	;
				14'b01001010111111: Data_out <= 16'h7B5F	;
				14'b01001011000000: Data_out <= 16'h7B5C	;
				14'b01001011000001: Data_out <= 16'h7B59	;
				14'b01001011000010: Data_out <= 16'h7B55	;
				14'b01001011000011: Data_out <= 16'h7B52	;
				14'b01001011000100: Data_out <= 16'h7B4F	;
				14'b01001011000101: Data_out <= 16'h7B4B	;
				14'b01001011000110: Data_out <= 16'h7B48	;
				14'b01001011000111: Data_out <= 16'h7B45	;
				14'b01001011001000: Data_out <= 16'h7B41	;
				14'b01001011001001: Data_out <= 16'h7B3E	;
				14'b01001011001010: Data_out <= 16'h7B3A	;
				14'b01001011001011: Data_out <= 16'h7B37	;
				14'b01001011001100: Data_out <= 16'h7B34	;
				14'b01001011001101: Data_out <= 16'h7B30	;
				14'b01001011001110: Data_out <= 16'h7B2D	;
				14'b01001011001111: Data_out <= 16'h7B29	;
				14'b01001011010000: Data_out <= 16'h7B26	;
				14'b01001011010001: Data_out <= 16'h7B23	;
				14'b01001011010010: Data_out <= 16'h7B1F	;
				14'b01001011010011: Data_out <= 16'h7B1C	;
				14'b01001011010100: Data_out <= 16'h7B18	;
				14'b01001011010101: Data_out <= 16'h7B15	;
				14'b01001011010110: Data_out <= 16'h7B11	;
				14'b01001011010111: Data_out <= 16'h7B0E	;
				14'b01001011011000: Data_out <= 16'h7B0A	;
				14'b01001011011001: Data_out <= 16'h7B07	;
				14'b01001011011010: Data_out <= 16'h7B03	;
				14'b01001011011011: Data_out <= 16'h7B00	;
				14'b01001011011100: Data_out <= 16'h7AFC	;
				14'b01001011011101: Data_out <= 16'h7AF9	;
				14'b01001011011110: Data_out <= 16'h7AF6	;
				14'b01001011011111: Data_out <= 16'h7AF2	;
				14'b01001011100000: Data_out <= 16'h7AEF	;
				14'b01001011100001: Data_out <= 16'h7AEB	;
				14'b01001011100010: Data_out <= 16'h7AE8	;
				14'b01001011100011: Data_out <= 16'h7AE4	;
				14'b01001011100100: Data_out <= 16'h7AE0	;
				14'b01001011100101: Data_out <= 16'h7ADD	;
				14'b01001011100110: Data_out <= 16'h7AD9	;
				14'b01001011100111: Data_out <= 16'h7AD6	;
				14'b01001011101000: Data_out <= 16'h7AD2	;
				14'b01001011101001: Data_out <= 16'h7ACF	;
				14'b01001011101010: Data_out <= 16'h7ACB	;
				14'b01001011101011: Data_out <= 16'h7AC8	;
				14'b01001011101100: Data_out <= 16'h7AC4	;
				14'b01001011101101: Data_out <= 16'h7AC1	;
				14'b01001011101110: Data_out <= 16'h7ABD	;
				14'b01001011101111: Data_out <= 16'h7ABA	;
				14'b01001011110000: Data_out <= 16'h7AB6	;
				14'b01001011110001: Data_out <= 16'h7AB2	;
				14'b01001011110010: Data_out <= 16'h7AAF	;
				14'b01001011110011: Data_out <= 16'h7AAB	;
				14'b01001011110100: Data_out <= 16'h7AA8	;
				14'b01001011110101: Data_out <= 16'h7AA4	;
				14'b01001011110110: Data_out <= 16'h7AA0	;
				14'b01001011110111: Data_out <= 16'h7A9D	;
				14'b01001011111000: Data_out <= 16'h7A99	;
				14'b01001011111001: Data_out <= 16'h7A96	;
				14'b01001011111010: Data_out <= 16'h7A92	;
				14'b01001011111011: Data_out <= 16'h7A8E	;
				14'b01001011111100: Data_out <= 16'h7A8B	;
				14'b01001011111101: Data_out <= 16'h7A87	;
				14'b01001011111110: Data_out <= 16'h7A83	;
				14'b01001011111111: Data_out <= 16'h7A80	;
				14'b01001100000000: Data_out <= 16'h7A7C	;
				14'b01001100000001: Data_out <= 16'h7A79	;
				14'b01001100000010: Data_out <= 16'h7A75	;
				14'b01001100000011: Data_out <= 16'h7A71	;
				14'b01001100000100: Data_out <= 16'h7A6E	;
				14'b01001100000101: Data_out <= 16'h7A6A	;
				14'b01001100000110: Data_out <= 16'h7A66	;
				14'b01001100000111: Data_out <= 16'h7A63	;
				14'b01001100001000: Data_out <= 16'h7A5F	;
				14'b01001100001001: Data_out <= 16'h7A5B	;
				14'b01001100001010: Data_out <= 16'h7A57	;
				14'b01001100001011: Data_out <= 16'h7A54	;
				14'b01001100001100: Data_out <= 16'h7A50	;
				14'b01001100001101: Data_out <= 16'h7A4C	;
				14'b01001100001110: Data_out <= 16'h7A49	;
				14'b01001100001111: Data_out <= 16'h7A45	;
				14'b01001100010000: Data_out <= 16'h7A41	;
				14'b01001100010001: Data_out <= 16'h7A3D	;
				14'b01001100010010: Data_out <= 16'h7A3A	;
				14'b01001100010011: Data_out <= 16'h7A36	;
				14'b01001100010100: Data_out <= 16'h7A32	;
				14'b01001100010101: Data_out <= 16'h7A2F	;
				14'b01001100010110: Data_out <= 16'h7A2B	;
				14'b01001100010111: Data_out <= 16'h7A27	;
				14'b01001100011000: Data_out <= 16'h7A23	;
				14'b01001100011001: Data_out <= 16'h7A20	;
				14'b01001100011010: Data_out <= 16'h7A1C	;
				14'b01001100011011: Data_out <= 16'h7A18	;
				14'b01001100011100: Data_out <= 16'h7A14	;
				14'b01001100011101: Data_out <= 16'h7A10	;
				14'b01001100011110: Data_out <= 16'h7A0D	;
				14'b01001100011111: Data_out <= 16'h7A09	;
				14'b01001100100000: Data_out <= 16'h7A05	;
				14'b01001100100001: Data_out <= 16'h7A01	;
				14'b01001100100010: Data_out <= 16'h79FD	;
				14'b01001100100011: Data_out <= 16'h79FA	;
				14'b01001100100100: Data_out <= 16'h79F6	;
				14'b01001100100101: Data_out <= 16'h79F2	;
				14'b01001100100110: Data_out <= 16'h79EE	;
				14'b01001100100111: Data_out <= 16'h79EA	;
				14'b01001100101000: Data_out <= 16'h79E7	;
				14'b01001100101001: Data_out <= 16'h79E3	;
				14'b01001100101010: Data_out <= 16'h79DF	;
				14'b01001100101011: Data_out <= 16'h79DB	;
				14'b01001100101100: Data_out <= 16'h79D7	;
				14'b01001100101101: Data_out <= 16'h79D3	;
				14'b01001100101110: Data_out <= 16'h79CF	;
				14'b01001100101111: Data_out <= 16'h79CC	;
				14'b01001100110000: Data_out <= 16'h79C8	;
				14'b01001100110001: Data_out <= 16'h79C4	;
				14'b01001100110010: Data_out <= 16'h79C0	;
				14'b01001100110011: Data_out <= 16'h79BC	;
				14'b01001100110100: Data_out <= 16'h79B8	;
				14'b01001100110101: Data_out <= 16'h79B4	;
				14'b01001100110110: Data_out <= 16'h79B0	;
				14'b01001100110111: Data_out <= 16'h79AD	;
				14'b01001100111000: Data_out <= 16'h79A9	;
				14'b01001100111001: Data_out <= 16'h79A5	;
				14'b01001100111010: Data_out <= 16'h79A1	;
				14'b01001100111011: Data_out <= 16'h799D	;
				14'b01001100111100: Data_out <= 16'h7999	;
				14'b01001100111101: Data_out <= 16'h7995	;
				14'b01001100111110: Data_out <= 16'h7991	;
				14'b01001100111111: Data_out <= 16'h798D	;
				14'b01001101000000: Data_out <= 16'h7989	;
				14'b01001101000001: Data_out <= 16'h7985	;
				14'b01001101000010: Data_out <= 16'h7981	;
				14'b01001101000011: Data_out <= 16'h797D	;
				14'b01001101000100: Data_out <= 16'h7979	;
				14'b01001101000101: Data_out <= 16'h7976	;
				14'b01001101000110: Data_out <= 16'h7972	;
				14'b01001101000111: Data_out <= 16'h796E	;
				14'b01001101001000: Data_out <= 16'h796A	;
				14'b01001101001001: Data_out <= 16'h7966	;
				14'b01001101001010: Data_out <= 16'h7962	;
				14'b01001101001011: Data_out <= 16'h795E	;
				14'b01001101001100: Data_out <= 16'h795A	;
				14'b01001101001101: Data_out <= 16'h7956	;
				14'b01001101001110: Data_out <= 16'h7952	;
				14'b01001101001111: Data_out <= 16'h794E	;
				14'b01001101010000: Data_out <= 16'h794A	;
				14'b01001101010001: Data_out <= 16'h7946	;
				14'b01001101010010: Data_out <= 16'h7942	;
				14'b01001101010011: Data_out <= 16'h793E	;
				14'b01001101010100: Data_out <= 16'h793A	;
				14'b01001101010101: Data_out <= 16'h7936	;
				14'b01001101010110: Data_out <= 16'h7931	;
				14'b01001101010111: Data_out <= 16'h792D	;
				14'b01001101011000: Data_out <= 16'h7929	;
				14'b01001101011001: Data_out <= 16'h7925	;
				14'b01001101011010: Data_out <= 16'h7921	;
				14'b01001101011011: Data_out <= 16'h791D	;
				14'b01001101011100: Data_out <= 16'h7919	;
				14'b01001101011101: Data_out <= 16'h7915	;
				14'b01001101011110: Data_out <= 16'h7911	;
				14'b01001101011111: Data_out <= 16'h790D	;
				14'b01001101100000: Data_out <= 16'h7909	;
				14'b01001101100001: Data_out <= 16'h7905	;
				14'b01001101100010: Data_out <= 16'h7901	;
				14'b01001101100011: Data_out <= 16'h78FD	;
				14'b01001101100100: Data_out <= 16'h78F8	;
				14'b01001101100101: Data_out <= 16'h78F4	;
				14'b01001101100110: Data_out <= 16'h78F0	;
				14'b01001101100111: Data_out <= 16'h78EC	;
				14'b01001101101000: Data_out <= 16'h78E8	;
				14'b01001101101001: Data_out <= 16'h78E4	;
				14'b01001101101010: Data_out <= 16'h78E0	;
				14'b01001101101011: Data_out <= 16'h78DC	;
				14'b01001101101100: Data_out <= 16'h78D7	;
				14'b01001101101101: Data_out <= 16'h78D3	;
				14'b01001101101110: Data_out <= 16'h78CF	;
				14'b01001101101111: Data_out <= 16'h78CB	;
				14'b01001101110000: Data_out <= 16'h78C7	;
				14'b01001101110001: Data_out <= 16'h78C3	;
				14'b01001101110010: Data_out <= 16'h78BE	;
				14'b01001101110011: Data_out <= 16'h78BA	;
				14'b01001101110100: Data_out <= 16'h78B6	;
				14'b01001101110101: Data_out <= 16'h78B2	;
				14'b01001101110110: Data_out <= 16'h78AE	;
				14'b01001101110111: Data_out <= 16'h78AA	;
				14'b01001101111000: Data_out <= 16'h78A5	;
				14'b01001101111001: Data_out <= 16'h78A1	;
				14'b01001101111010: Data_out <= 16'h789D	;
				14'b01001101111011: Data_out <= 16'h7899	;
				14'b01001101111100: Data_out <= 16'h7895	;
				14'b01001101111101: Data_out <= 16'h7890	;
				14'b01001101111110: Data_out <= 16'h788C	;
				14'b01001101111111: Data_out <= 16'h7888	;
				14'b01001110000000: Data_out <= 16'h7884	;
				14'b01001110000001: Data_out <= 16'h787F	;
				14'b01001110000010: Data_out <= 16'h787B	;
				14'b01001110000011: Data_out <= 16'h7877	;
				14'b01001110000100: Data_out <= 16'h7873	;
				14'b01001110000101: Data_out <= 16'h786E	;
				14'b01001110000110: Data_out <= 16'h786A	;
				14'b01001110000111: Data_out <= 16'h7866	;
				14'b01001110001000: Data_out <= 16'h7862	;
				14'b01001110001001: Data_out <= 16'h785D	;
				14'b01001110001010: Data_out <= 16'h7859	;
				14'b01001110001011: Data_out <= 16'h7855	;
				14'b01001110001100: Data_out <= 16'h7851	;
				14'b01001110001101: Data_out <= 16'h784C	;
				14'b01001110001110: Data_out <= 16'h7848	;
				14'b01001110001111: Data_out <= 16'h7844	;
				14'b01001110010000: Data_out <= 16'h783F	;
				14'b01001110010001: Data_out <= 16'h783B	;
				14'b01001110010010: Data_out <= 16'h7837	;
				14'b01001110010011: Data_out <= 16'h7832	;
				14'b01001110010100: Data_out <= 16'h782E	;
				14'b01001110010101: Data_out <= 16'h782A	;
				14'b01001110010110: Data_out <= 16'h7825	;
				14'b01001110010111: Data_out <= 16'h7821	;
				14'b01001110011000: Data_out <= 16'h781D	;
				14'b01001110011001: Data_out <= 16'h7818	;
				14'b01001110011010: Data_out <= 16'h7814	;
				14'b01001110011011: Data_out <= 16'h7810	;
				14'b01001110011100: Data_out <= 16'h780B	;
				14'b01001110011101: Data_out <= 16'h7807	;
				14'b01001110011110: Data_out <= 16'h7803	;
				14'b01001110011111: Data_out <= 16'h77FE	;
				14'b01001110100000: Data_out <= 16'h77FA	;
				14'b01001110100001: Data_out <= 16'h77F6	;
				14'b01001110100010: Data_out <= 16'h77F1	;
				14'b01001110100011: Data_out <= 16'h77ED	;
				14'b01001110100100: Data_out <= 16'h77E8	;
				14'b01001110100101: Data_out <= 16'h77E4	;
				14'b01001110100110: Data_out <= 16'h77E0	;
				14'b01001110100111: Data_out <= 16'h77DB	;
				14'b01001110101000: Data_out <= 16'h77D7	;
				14'b01001110101001: Data_out <= 16'h77D2	;
				14'b01001110101010: Data_out <= 16'h77CE	;
				14'b01001110101011: Data_out <= 16'h77C9	;
				14'b01001110101100: Data_out <= 16'h77C5	;
				14'b01001110101101: Data_out <= 16'h77C1	;
				14'b01001110101110: Data_out <= 16'h77BC	;
				14'b01001110101111: Data_out <= 16'h77B8	;
				14'b01001110110000: Data_out <= 16'h77B3	;
				14'b01001110110001: Data_out <= 16'h77AF	;
				14'b01001110110010: Data_out <= 16'h77AA	;
				14'b01001110110011: Data_out <= 16'h77A6	;
				14'b01001110110100: Data_out <= 16'h77A1	;
				14'b01001110110101: Data_out <= 16'h779D	;
				14'b01001110110110: Data_out <= 16'h7798	;
				14'b01001110110111: Data_out <= 16'h7794	;
				14'b01001110111000: Data_out <= 16'h7790	;
				14'b01001110111001: Data_out <= 16'h778B	;
				14'b01001110111010: Data_out <= 16'h7787	;
				14'b01001110111011: Data_out <= 16'h7782	;
				14'b01001110111100: Data_out <= 16'h777E	;
				14'b01001110111101: Data_out <= 16'h7779	;
				14'b01001110111110: Data_out <= 16'h7775	;
				14'b01001110111111: Data_out <= 16'h7770	;
				14'b01001111000000: Data_out <= 16'h776B	;
				14'b01001111000001: Data_out <= 16'h7767	;
				14'b01001111000010: Data_out <= 16'h7762	;
				14'b01001111000011: Data_out <= 16'h775E	;
				14'b01001111000100: Data_out <= 16'h7759	;
				14'b01001111000101: Data_out <= 16'h7755	;
				14'b01001111000110: Data_out <= 16'h7750	;
				14'b01001111000111: Data_out <= 16'h774C	;
				14'b01001111001000: Data_out <= 16'h7747	;
				14'b01001111001001: Data_out <= 16'h7743	;
				14'b01001111001010: Data_out <= 16'h773E	;
				14'b01001111001011: Data_out <= 16'h7739	;
				14'b01001111001100: Data_out <= 16'h7735	;
				14'b01001111001101: Data_out <= 16'h7730	;
				14'b01001111001110: Data_out <= 16'h772C	;
				14'b01001111001111: Data_out <= 16'h7727	;
				14'b01001111010000: Data_out <= 16'h7723	;
				14'b01001111010001: Data_out <= 16'h771E	;
				14'b01001111010010: Data_out <= 16'h7719	;
				14'b01001111010011: Data_out <= 16'h7715	;
				14'b01001111010100: Data_out <= 16'h7710	;
				14'b01001111010101: Data_out <= 16'h770C	;
				14'b01001111010110: Data_out <= 16'h7707	;
				14'b01001111010111: Data_out <= 16'h7702	;
				14'b01001111011000: Data_out <= 16'h76FE	;
				14'b01001111011001: Data_out <= 16'h76F9	;
				14'b01001111011010: Data_out <= 16'h76F4	;
				14'b01001111011011: Data_out <= 16'h76F0	;
				14'b01001111011100: Data_out <= 16'h76EB	;
				14'b01001111011101: Data_out <= 16'h76E6	;
				14'b01001111011110: Data_out <= 16'h76E2	;
				14'b01001111011111: Data_out <= 16'h76DD	;
				14'b01001111100000: Data_out <= 16'h76D8	;
				14'b01001111100001: Data_out <= 16'h76D4	;
				14'b01001111100010: Data_out <= 16'h76CF	;
				14'b01001111100011: Data_out <= 16'h76CA	;
				14'b01001111100100: Data_out <= 16'h76C6	;
				14'b01001111100101: Data_out <= 16'h76C1	;
				14'b01001111100110: Data_out <= 16'h76BC	;
				14'b01001111100111: Data_out <= 16'h76B8	;
				14'b01001111101000: Data_out <= 16'h76B3	;
				14'b01001111101001: Data_out <= 16'h76AE	;
				14'b01001111101010: Data_out <= 16'h76AA	;
				14'b01001111101011: Data_out <= 16'h76A5	;
				14'b01001111101100: Data_out <= 16'h76A0	;
				14'b01001111101101: Data_out <= 16'h769B	;
				14'b01001111101110: Data_out <= 16'h7697	;
				14'b01001111101111: Data_out <= 16'h7692	;
				14'b01001111110000: Data_out <= 16'h768D	;
				14'b01001111110001: Data_out <= 16'h7688	;
				14'b01001111110010: Data_out <= 16'h7684	;
				14'b01001111110011: Data_out <= 16'h767F	;
				14'b01001111110100: Data_out <= 16'h767A	;
				14'b01001111110101: Data_out <= 16'h7675	;
				14'b01001111110110: Data_out <= 16'h7671	;
				14'b01001111110111: Data_out <= 16'h766C	;
				14'b01001111111000: Data_out <= 16'h7667	;
				14'b01001111111001: Data_out <= 16'h7662	;
				14'b01001111111010: Data_out <= 16'h765E	;
				14'b01001111111011: Data_out <= 16'h7659	;
				14'b01001111111100: Data_out <= 16'h7654	;
				14'b01001111111101: Data_out <= 16'h764F	;
				14'b01001111111110: Data_out <= 16'h764A	;
				14'b01001111111111: Data_out <= 16'h7646	;
				14'b01010000000000: Data_out <= 16'h7641	;
				14'b01010000000001: Data_out <= 16'h763C	;
				14'b01010000000010: Data_out <= 16'h7637	;
				14'b01010000000011: Data_out <= 16'h7632	;
				14'b01010000000100: Data_out <= 16'h762E	;
				14'b01010000000101: Data_out <= 16'h7629	;
				14'b01010000000110: Data_out <= 16'h7624	;
				14'b01010000000111: Data_out <= 16'h761F	;
				14'b01010000001000: Data_out <= 16'h761A	;
				14'b01010000001001: Data_out <= 16'h7615	;
				14'b01010000001010: Data_out <= 16'h7611	;
				14'b01010000001011: Data_out <= 16'h760C	;
				14'b01010000001100: Data_out <= 16'h7607	;
				14'b01010000001101: Data_out <= 16'h7602	;
				14'b01010000001110: Data_out <= 16'h75FD	;
				14'b01010000001111: Data_out <= 16'h75F8	;
				14'b01010000010000: Data_out <= 16'h75F3	;
				14'b01010000010001: Data_out <= 16'h75EE	;
				14'b01010000010010: Data_out <= 16'h75EA	;
				14'b01010000010011: Data_out <= 16'h75E5	;
				14'b01010000010100: Data_out <= 16'h75E0	;
				14'b01010000010101: Data_out <= 16'h75DB	;
				14'b01010000010110: Data_out <= 16'h75D6	;
				14'b01010000010111: Data_out <= 16'h75D1	;
				14'b01010000011000: Data_out <= 16'h75CC	;
				14'b01010000011001: Data_out <= 16'h75C7	;
				14'b01010000011010: Data_out <= 16'h75C2	;
				14'b01010000011011: Data_out <= 16'h75BD	;
				14'b01010000011100: Data_out <= 16'h75B8	;
				14'b01010000011101: Data_out <= 16'h75B4	;
				14'b01010000011110: Data_out <= 16'h75AF	;
				14'b01010000011111: Data_out <= 16'h75AA	;
				14'b01010000100000: Data_out <= 16'h75A5	;
				14'b01010000100001: Data_out <= 16'h75A0	;
				14'b01010000100010: Data_out <= 16'h759B	;
				14'b01010000100011: Data_out <= 16'h7596	;
				14'b01010000100100: Data_out <= 16'h7591	;
				14'b01010000100101: Data_out <= 16'h758C	;
				14'b01010000100110: Data_out <= 16'h7587	;
				14'b01010000100111: Data_out <= 16'h7582	;
				14'b01010000101000: Data_out <= 16'h757D	;
				14'b01010000101001: Data_out <= 16'h7578	;
				14'b01010000101010: Data_out <= 16'h7573	;
				14'b01010000101011: Data_out <= 16'h756E	;
				14'b01010000101100: Data_out <= 16'h7569	;
				14'b01010000101101: Data_out <= 16'h7564	;
				14'b01010000101110: Data_out <= 16'h755F	;
				14'b01010000101111: Data_out <= 16'h755A	;
				14'b01010000110000: Data_out <= 16'h7555	;
				14'b01010000110001: Data_out <= 16'h7550	;
				14'b01010000110010: Data_out <= 16'h754B	;
				14'b01010000110011: Data_out <= 16'h7546	;
				14'b01010000110100: Data_out <= 16'h7541	;
				14'b01010000110101: Data_out <= 16'h753C	;
				14'b01010000110110: Data_out <= 16'h7537	;
				14'b01010000110111: Data_out <= 16'h7532	;
				14'b01010000111000: Data_out <= 16'h752D	;
				14'b01010000111001: Data_out <= 16'h7528	;
				14'b01010000111010: Data_out <= 16'h7522	;
				14'b01010000111011: Data_out <= 16'h751D	;
				14'b01010000111100: Data_out <= 16'h7518	;
				14'b01010000111101: Data_out <= 16'h7513	;
				14'b01010000111110: Data_out <= 16'h750E	;
				14'b01010000111111: Data_out <= 16'h7509	;
				14'b01010001000000: Data_out <= 16'h7504	;
				14'b01010001000001: Data_out <= 16'h74FF	;
				14'b01010001000010: Data_out <= 16'h74FA	;
				14'b01010001000011: Data_out <= 16'h74F5	;
				14'b01010001000100: Data_out <= 16'h74F0	;
				14'b01010001000101: Data_out <= 16'h74EA	;
				14'b01010001000110: Data_out <= 16'h74E5	;
				14'b01010001000111: Data_out <= 16'h74E0	;
				14'b01010001001000: Data_out <= 16'h74DB	;
				14'b01010001001001: Data_out <= 16'h74D6	;
				14'b01010001001010: Data_out <= 16'h74D1	;
				14'b01010001001011: Data_out <= 16'h74CC	;
				14'b01010001001100: Data_out <= 16'h74C7	;
				14'b01010001001101: Data_out <= 16'h74C1	;
				14'b01010001001110: Data_out <= 16'h74BC	;
				14'b01010001001111: Data_out <= 16'h74B7	;
				14'b01010001010000: Data_out <= 16'h74B2	;
				14'b01010001010001: Data_out <= 16'h74AD	;
				14'b01010001010010: Data_out <= 16'h74A8	;
				14'b01010001010011: Data_out <= 16'h74A2	;
				14'b01010001010100: Data_out <= 16'h749D	;
				14'b01010001010101: Data_out <= 16'h7498	;
				14'b01010001010110: Data_out <= 16'h7493	;
				14'b01010001010111: Data_out <= 16'h748E	;
				14'b01010001011000: Data_out <= 16'h7489	;
				14'b01010001011001: Data_out <= 16'h7483	;
				14'b01010001011010: Data_out <= 16'h747E	;
				14'b01010001011011: Data_out <= 16'h7479	;
				14'b01010001011100: Data_out <= 16'h7474	;
				14'b01010001011101: Data_out <= 16'h746E	;
				14'b01010001011110: Data_out <= 16'h7469	;
				14'b01010001011111: Data_out <= 16'h7464	;
				14'b01010001100000: Data_out <= 16'h745F	;
				14'b01010001100001: Data_out <= 16'h745A	;
				14'b01010001100010: Data_out <= 16'h7454	;
				14'b01010001100011: Data_out <= 16'h744F	;
				14'b01010001100100: Data_out <= 16'h744A	;
				14'b01010001100101: Data_out <= 16'h7445	;
				14'b01010001100110: Data_out <= 16'h743F	;
				14'b01010001100111: Data_out <= 16'h743A	;
				14'b01010001101000: Data_out <= 16'h7435	;
				14'b01010001101001: Data_out <= 16'h7430	;
				14'b01010001101010: Data_out <= 16'h742A	;
				14'b01010001101011: Data_out <= 16'h7425	;
				14'b01010001101100: Data_out <= 16'h7420	;
				14'b01010001101101: Data_out <= 16'h741A	;
				14'b01010001101110: Data_out <= 16'h7415	;
				14'b01010001101111: Data_out <= 16'h7410	;
				14'b01010001110000: Data_out <= 16'h740B	;
				14'b01010001110001: Data_out <= 16'h7405	;
				14'b01010001110010: Data_out <= 16'h7400	;
				14'b01010001110011: Data_out <= 16'h73FB	;
				14'b01010001110100: Data_out <= 16'h73F5	;
				14'b01010001110101: Data_out <= 16'h73F0	;
				14'b01010001110110: Data_out <= 16'h73EB	;
				14'b01010001110111: Data_out <= 16'h73E5	;
				14'b01010001111000: Data_out <= 16'h73E0	;
				14'b01010001111001: Data_out <= 16'h73DB	;
				14'b01010001111010: Data_out <= 16'h73D5	;
				14'b01010001111011: Data_out <= 16'h73D0	;
				14'b01010001111100: Data_out <= 16'h73CB	;
				14'b01010001111101: Data_out <= 16'h73C5	;
				14'b01010001111110: Data_out <= 16'h73C0	;
				14'b01010001111111: Data_out <= 16'h73BA	;
				14'b01010010000000: Data_out <= 16'h73B5	;
				14'b01010010000001: Data_out <= 16'h73B0	;
				14'b01010010000010: Data_out <= 16'h73AA	;
				14'b01010010000011: Data_out <= 16'h73A5	;
				14'b01010010000100: Data_out <= 16'h73A0	;
				14'b01010010000101: Data_out <= 16'h739A	;
				14'b01010010000110: Data_out <= 16'h7395	;
				14'b01010010000111: Data_out <= 16'h738F	;
				14'b01010010001000: Data_out <= 16'h738A	;
				14'b01010010001001: Data_out <= 16'h7385	;
				14'b01010010001010: Data_out <= 16'h737F	;
				14'b01010010001011: Data_out <= 16'h737A	;
				14'b01010010001100: Data_out <= 16'h7374	;
				14'b01010010001101: Data_out <= 16'h736F	;
				14'b01010010001110: Data_out <= 16'h7369	;
				14'b01010010001111: Data_out <= 16'h7364	;
				14'b01010010010000: Data_out <= 16'h735F	;
				14'b01010010010001: Data_out <= 16'h7359	;
				14'b01010010010010: Data_out <= 16'h7354	;
				14'b01010010010011: Data_out <= 16'h734E	;
				14'b01010010010100: Data_out <= 16'h7349	;
				14'b01010010010101: Data_out <= 16'h7343	;
				14'b01010010010110: Data_out <= 16'h733E	;
				14'b01010010010111: Data_out <= 16'h7338	;
				14'b01010010011000: Data_out <= 16'h7333	;
				14'b01010010011001: Data_out <= 16'h732D	;
				14'b01010010011010: Data_out <= 16'h7328	;
				14'b01010010011011: Data_out <= 16'h7322	;
				14'b01010010011100: Data_out <= 16'h731D	;
				14'b01010010011101: Data_out <= 16'h7317	;
				14'b01010010011110: Data_out <= 16'h7312	;
				14'b01010010011111: Data_out <= 16'h730C	;
				14'b01010010100000: Data_out <= 16'h7307	;
				14'b01010010100001: Data_out <= 16'h7301	;
				14'b01010010100010: Data_out <= 16'h72FC	;
				14'b01010010100011: Data_out <= 16'h72F6	;
				14'b01010010100100: Data_out <= 16'h72F1	;
				14'b01010010100101: Data_out <= 16'h72EB	;
				14'b01010010100110: Data_out <= 16'h72E6	;
				14'b01010010100111: Data_out <= 16'h72E0	;
				14'b01010010101000: Data_out <= 16'h72DB	;
				14'b01010010101001: Data_out <= 16'h72D5	;
				14'b01010010101010: Data_out <= 16'h72D0	;
				14'b01010010101011: Data_out <= 16'h72CA	;
				14'b01010010101100: Data_out <= 16'h72C5	;
				14'b01010010101101: Data_out <= 16'h72BF	;
				14'b01010010101110: Data_out <= 16'h72B9	;
				14'b01010010101111: Data_out <= 16'h72B4	;
				14'b01010010110000: Data_out <= 16'h72AE	;
				14'b01010010110001: Data_out <= 16'h72A9	;
				14'b01010010110010: Data_out <= 16'h72A3	;
				14'b01010010110011: Data_out <= 16'h729D	;
				14'b01010010110100: Data_out <= 16'h7298	;
				14'b01010010110101: Data_out <= 16'h7292	;
				14'b01010010110110: Data_out <= 16'h728D	;
				14'b01010010110111: Data_out <= 16'h7287	;
				14'b01010010111000: Data_out <= 16'h7281	;
				14'b01010010111001: Data_out <= 16'h727C	;
				14'b01010010111010: Data_out <= 16'h7276	;
				14'b01010010111011: Data_out <= 16'h7271	;
				14'b01010010111100: Data_out <= 16'h726B	;
				14'b01010010111101: Data_out <= 16'h7265	;
				14'b01010010111110: Data_out <= 16'h7260	;
				14'b01010010111111: Data_out <= 16'h725A	;
				14'b01010011000000: Data_out <= 16'h7254	;
				14'b01010011000001: Data_out <= 16'h724F	;
				14'b01010011000010: Data_out <= 16'h7249	;
				14'b01010011000011: Data_out <= 16'h7243	;
				14'b01010011000100: Data_out <= 16'h723E	;
				14'b01010011000101: Data_out <= 16'h7238	;
				14'b01010011000110: Data_out <= 16'h7232	;
				14'b01010011000111: Data_out <= 16'h722D	;
				14'b01010011001000: Data_out <= 16'h7227	;
				14'b01010011001001: Data_out <= 16'h7221	;
				14'b01010011001010: Data_out <= 16'h721C	;
				14'b01010011001011: Data_out <= 16'h7216	;
				14'b01010011001100: Data_out <= 16'h7210	;
				14'b01010011001101: Data_out <= 16'h720B	;
				14'b01010011001110: Data_out <= 16'h7205	;
				14'b01010011001111: Data_out <= 16'h71FF	;
				14'b01010011010000: Data_out <= 16'h71F9	;
				14'b01010011010001: Data_out <= 16'h71F4	;
				14'b01010011010010: Data_out <= 16'h71EE	;
				14'b01010011010011: Data_out <= 16'h71E8	;
				14'b01010011010100: Data_out <= 16'h71E3	;
				14'b01010011010101: Data_out <= 16'h71DD	;
				14'b01010011010110: Data_out <= 16'h71D7	;
				14'b01010011010111: Data_out <= 16'h71D1	;
				14'b01010011011000: Data_out <= 16'h71CC	;
				14'b01010011011001: Data_out <= 16'h71C6	;
				14'b01010011011010: Data_out <= 16'h71C0	;
				14'b01010011011011: Data_out <= 16'h71BA	;
				14'b01010011011100: Data_out <= 16'h71B5	;
				14'b01010011011101: Data_out <= 16'h71AF	;
				14'b01010011011110: Data_out <= 16'h71A9	;
				14'b01010011011111: Data_out <= 16'h71A3	;
				14'b01010011100000: Data_out <= 16'h719D	;
				14'b01010011100001: Data_out <= 16'h7198	;
				14'b01010011100010: Data_out <= 16'h7192	;
				14'b01010011100011: Data_out <= 16'h718C	;
				14'b01010011100100: Data_out <= 16'h7186	;
				14'b01010011100101: Data_out <= 16'h7180	;
				14'b01010011100110: Data_out <= 16'h717B	;
				14'b01010011100111: Data_out <= 16'h7175	;
				14'b01010011101000: Data_out <= 16'h716F	;
				14'b01010011101001: Data_out <= 16'h7169	;
				14'b01010011101010: Data_out <= 16'h7163	;
				14'b01010011101011: Data_out <= 16'h715D	;
				14'b01010011101100: Data_out <= 16'h7158	;
				14'b01010011101101: Data_out <= 16'h7152	;
				14'b01010011101110: Data_out <= 16'h714C	;
				14'b01010011101111: Data_out <= 16'h7146	;
				14'b01010011110000: Data_out <= 16'h7140	;
				14'b01010011110001: Data_out <= 16'h713A	;
				14'b01010011110010: Data_out <= 16'h7135	;
				14'b01010011110011: Data_out <= 16'h712F	;
				14'b01010011110100: Data_out <= 16'h7129	;
				14'b01010011110101: Data_out <= 16'h7123	;
				14'b01010011110110: Data_out <= 16'h711D	;
				14'b01010011110111: Data_out <= 16'h7117	;
				14'b01010011111000: Data_out <= 16'h7111	;
				14'b01010011111001: Data_out <= 16'h710B	;
				14'b01010011111010: Data_out <= 16'h7105	;
				14'b01010011111011: Data_out <= 16'h7100	;
				14'b01010011111100: Data_out <= 16'h70FA	;
				14'b01010011111101: Data_out <= 16'h70F4	;
				14'b01010011111110: Data_out <= 16'h70EE	;
				14'b01010011111111: Data_out <= 16'h70E8	;
				14'b01010100000000: Data_out <= 16'h70E2	;
				14'b01010100000001: Data_out <= 16'h70DC	;
				14'b01010100000010: Data_out <= 16'h70D6	;
				14'b01010100000011: Data_out <= 16'h70D0	;
				14'b01010100000100: Data_out <= 16'h70CA	;
				14'b01010100000101: Data_out <= 16'h70C4	;
				14'b01010100000110: Data_out <= 16'h70BE	;
				14'b01010100000111: Data_out <= 16'h70B8	;
				14'b01010100001000: Data_out <= 16'h70B2	;
				14'b01010100001001: Data_out <= 16'h70AD	;
				14'b01010100001010: Data_out <= 16'h70A7	;
				14'b01010100001011: Data_out <= 16'h70A1	;
				14'b01010100001100: Data_out <= 16'h709B	;
				14'b01010100001101: Data_out <= 16'h7095	;
				14'b01010100001110: Data_out <= 16'h708F	;
				14'b01010100001111: Data_out <= 16'h7089	;
				14'b01010100010000: Data_out <= 16'h7083	;
				14'b01010100010001: Data_out <= 16'h707D	;
				14'b01010100010010: Data_out <= 16'h7077	;
				14'b01010100010011: Data_out <= 16'h7071	;
				14'b01010100010100: Data_out <= 16'h706B	;
				14'b01010100010101: Data_out <= 16'h7065	;
				14'b01010100010110: Data_out <= 16'h705F	;
				14'b01010100010111: Data_out <= 16'h7059	;
				14'b01010100011000: Data_out <= 16'h7053	;
				14'b01010100011001: Data_out <= 16'h704D	;
				14'b01010100011010: Data_out <= 16'h7047	;
				14'b01010100011011: Data_out <= 16'h7041	;
				14'b01010100011100: Data_out <= 16'h703A	;
				14'b01010100011101: Data_out <= 16'h7034	;
				14'b01010100011110: Data_out <= 16'h702E	;
				14'b01010100011111: Data_out <= 16'h7028	;
				14'b01010100100000: Data_out <= 16'h7022	;
				14'b01010100100001: Data_out <= 16'h701C	;
				14'b01010100100010: Data_out <= 16'h7016	;
				14'b01010100100011: Data_out <= 16'h7010	;
				14'b01010100100100: Data_out <= 16'h700A	;
				14'b01010100100101: Data_out <= 16'h7004	;
				14'b01010100100110: Data_out <= 16'h6FFE	;
				14'b01010100100111: Data_out <= 16'h6FF8	;
				14'b01010100101000: Data_out <= 16'h6FF2	;
				14'b01010100101001: Data_out <= 16'h6FEC	;
				14'b01010100101010: Data_out <= 16'h6FE5	;
				14'b01010100101011: Data_out <= 16'h6FDF	;
				14'b01010100101100: Data_out <= 16'h6FD9	;
				14'b01010100101101: Data_out <= 16'h6FD3	;
				14'b01010100101110: Data_out <= 16'h6FCD	;
				14'b01010100101111: Data_out <= 16'h6FC7	;
				14'b01010100110000: Data_out <= 16'h6FC1	;
				14'b01010100110001: Data_out <= 16'h6FBB	;
				14'b01010100110010: Data_out <= 16'h6FB5	;
				14'b01010100110011: Data_out <= 16'h6FAE	;
				14'b01010100110100: Data_out <= 16'h6FA8	;
				14'b01010100110101: Data_out <= 16'h6FA2	;
				14'b01010100110110: Data_out <= 16'h6F9C	;
				14'b01010100110111: Data_out <= 16'h6F96	;
				14'b01010100111000: Data_out <= 16'h6F90	;
				14'b01010100111001: Data_out <= 16'h6F89	;
				14'b01010100111010: Data_out <= 16'h6F83	;
				14'b01010100111011: Data_out <= 16'h6F7D	;
				14'b01010100111100: Data_out <= 16'h6F77	;
				14'b01010100111101: Data_out <= 16'h6F71	;
				14'b01010100111110: Data_out <= 16'h6F6B	;
				14'b01010100111111: Data_out <= 16'h6F64	;
				14'b01010101000000: Data_out <= 16'h6F5E	;
				14'b01010101000001: Data_out <= 16'h6F58	;
				14'b01010101000010: Data_out <= 16'h6F52	;
				14'b01010101000011: Data_out <= 16'h6F4C	;
				14'b01010101000100: Data_out <= 16'h6F45	;
				14'b01010101000101: Data_out <= 16'h6F3F	;
				14'b01010101000110: Data_out <= 16'h6F39	;
				14'b01010101000111: Data_out <= 16'h6F33	;
				14'b01010101001000: Data_out <= 16'h6F2D	;
				14'b01010101001001: Data_out <= 16'h6F26	;
				14'b01010101001010: Data_out <= 16'h6F20	;
				14'b01010101001011: Data_out <= 16'h6F1A	;
				14'b01010101001100: Data_out <= 16'h6F14	;
				14'b01010101001101: Data_out <= 16'h6F0D	;
				14'b01010101001110: Data_out <= 16'h6F07	;
				14'b01010101001111: Data_out <= 16'h6F01	;
				14'b01010101010000: Data_out <= 16'h6EFB	;
				14'b01010101010001: Data_out <= 16'h6EF4	;
				14'b01010101010010: Data_out <= 16'h6EEE	;
				14'b01010101010011: Data_out <= 16'h6EE8	;
				14'b01010101010100: Data_out <= 16'h6EE2	;
				14'b01010101010101: Data_out <= 16'h6EDB	;
				14'b01010101010110: Data_out <= 16'h6ED5	;
				14'b01010101010111: Data_out <= 16'h6ECF	;
				14'b01010101011000: Data_out <= 16'h6EC8	;
				14'b01010101011001: Data_out <= 16'h6EC2	;
				14'b01010101011010: Data_out <= 16'h6EBC	;
				14'b01010101011011: Data_out <= 16'h6EB5	;
				14'b01010101011100: Data_out <= 16'h6EAF	;
				14'b01010101011101: Data_out <= 16'h6EA9	;
				14'b01010101011110: Data_out <= 16'h6EA3	;
				14'b01010101011111: Data_out <= 16'h6E9C	;
				14'b01010101100000: Data_out <= 16'h6E96	;
				14'b01010101100001: Data_out <= 16'h6E90	;
				14'b01010101100010: Data_out <= 16'h6E89	;
				14'b01010101100011: Data_out <= 16'h6E83	;
				14'b01010101100100: Data_out <= 16'h6E7D	;
				14'b01010101100101: Data_out <= 16'h6E76	;
				14'b01010101100110: Data_out <= 16'h6E70	;
				14'b01010101100111: Data_out <= 16'h6E6A	;
				14'b01010101101000: Data_out <= 16'h6E63	;
				14'b01010101101001: Data_out <= 16'h6E5D	;
				14'b01010101101010: Data_out <= 16'h6E56	;
				14'b01010101101011: Data_out <= 16'h6E50	;
				14'b01010101101100: Data_out <= 16'h6E4A	;
				14'b01010101101101: Data_out <= 16'h6E43	;
				14'b01010101101110: Data_out <= 16'h6E3D	;
				14'b01010101101111: Data_out <= 16'h6E37	;
				14'b01010101110000: Data_out <= 16'h6E30	;
				14'b01010101110001: Data_out <= 16'h6E2A	;
				14'b01010101110010: Data_out <= 16'h6E23	;
				14'b01010101110011: Data_out <= 16'h6E1D	;
				14'b01010101110100: Data_out <= 16'h6E17	;
				14'b01010101110101: Data_out <= 16'h6E10	;
				14'b01010101110110: Data_out <= 16'h6E0A	;
				14'b01010101110111: Data_out <= 16'h6E03	;
				14'b01010101111000: Data_out <= 16'h6DFD	;
				14'b01010101111001: Data_out <= 16'h6DF6	;
				14'b01010101111010: Data_out <= 16'h6DF0	;
				14'b01010101111011: Data_out <= 16'h6DEA	;
				14'b01010101111100: Data_out <= 16'h6DE3	;
				14'b01010101111101: Data_out <= 16'h6DDD	;
				14'b01010101111110: Data_out <= 16'h6DD6	;
				14'b01010101111111: Data_out <= 16'h6DD0	;
				14'b01010110000000: Data_out <= 16'h6DC9	;
				14'b01010110000001: Data_out <= 16'h6DC3	;
				14'b01010110000010: Data_out <= 16'h6DBC	;
				14'b01010110000011: Data_out <= 16'h6DB6	;
				14'b01010110000100: Data_out <= 16'h6DAF	;
				14'b01010110000101: Data_out <= 16'h6DA9	;
				14'b01010110000110: Data_out <= 16'h6DA2	;
				14'b01010110000111: Data_out <= 16'h6D9C	;
				14'b01010110001000: Data_out <= 16'h6D95	;
				14'b01010110001001: Data_out <= 16'h6D8F	;
				14'b01010110001010: Data_out <= 16'h6D88	;
				14'b01010110001011: Data_out <= 16'h6D82	;
				14'b01010110001100: Data_out <= 16'h6D7B	;
				14'b01010110001101: Data_out <= 16'h6D75	;
				14'b01010110001110: Data_out <= 16'h6D6E	;
				14'b01010110001111: Data_out <= 16'h6D68	;
				14'b01010110010000: Data_out <= 16'h6D61	;
				14'b01010110010001: Data_out <= 16'h6D5B	;
				14'b01010110010010: Data_out <= 16'h6D54	;
				14'b01010110010011: Data_out <= 16'h6D4E	;
				14'b01010110010100: Data_out <= 16'h6D47	;
				14'b01010110010101: Data_out <= 16'h6D41	;
				14'b01010110010110: Data_out <= 16'h6D3A	;
				14'b01010110010111: Data_out <= 16'h6D34	;
				14'b01010110011000: Data_out <= 16'h6D2D	;
				14'b01010110011001: Data_out <= 16'h6D26	;
				14'b01010110011010: Data_out <= 16'h6D20	;
				14'b01010110011011: Data_out <= 16'h6D19	;
				14'b01010110011100: Data_out <= 16'h6D13	;
				14'b01010110011101: Data_out <= 16'h6D0C	;
				14'b01010110011110: Data_out <= 16'h6D06	;
				14'b01010110011111: Data_out <= 16'h6CFF	;
				14'b01010110100000: Data_out <= 16'h6CF8	;
				14'b01010110100001: Data_out <= 16'h6CF2	;
				14'b01010110100010: Data_out <= 16'h6CEB	;
				14'b01010110100011: Data_out <= 16'h6CE5	;
				14'b01010110100100: Data_out <= 16'h6CDE	;
				14'b01010110100101: Data_out <= 16'h6CD7	;
				14'b01010110100110: Data_out <= 16'h6CD1	;
				14'b01010110100111: Data_out <= 16'h6CCA	;
				14'b01010110101000: Data_out <= 16'h6CC4	;
				14'b01010110101001: Data_out <= 16'h6CBD	;
				14'b01010110101010: Data_out <= 16'h6CB6	;
				14'b01010110101011: Data_out <= 16'h6CB0	;
				14'b01010110101100: Data_out <= 16'h6CA9	;
				14'b01010110101101: Data_out <= 16'h6CA2	;
				14'b01010110101110: Data_out <= 16'h6C9C	;
				14'b01010110101111: Data_out <= 16'h6C95	;
				14'b01010110110000: Data_out <= 16'h6C8E	;
				14'b01010110110001: Data_out <= 16'h6C88	;
				14'b01010110110010: Data_out <= 16'h6C81	;
				14'b01010110110011: Data_out <= 16'h6C7A	;
				14'b01010110110100: Data_out <= 16'h6C74	;
				14'b01010110110101: Data_out <= 16'h6C6D	;
				14'b01010110110110: Data_out <= 16'h6C66	;
				14'b01010110110111: Data_out <= 16'h6C60	;
				14'b01010110111000: Data_out <= 16'h6C59	;
				14'b01010110111001: Data_out <= 16'h6C52	;
				14'b01010110111010: Data_out <= 16'h6C4C	;
				14'b01010110111011: Data_out <= 16'h6C45	;
				14'b01010110111100: Data_out <= 16'h6C3E	;
				14'b01010110111101: Data_out <= 16'h6C38	;
				14'b01010110111110: Data_out <= 16'h6C31	;
				14'b01010110111111: Data_out <= 16'h6C2A	;
				14'b01010111000000: Data_out <= 16'h6C23	;
				14'b01010111000001: Data_out <= 16'h6C1D	;
				14'b01010111000010: Data_out <= 16'h6C16	;
				14'b01010111000011: Data_out <= 16'h6C0F	;
				14'b01010111000100: Data_out <= 16'h6C08	;
				14'b01010111000101: Data_out <= 16'h6C02	;
				14'b01010111000110: Data_out <= 16'h6BFB	;
				14'b01010111000111: Data_out <= 16'h6BF4	;
				14'b01010111001000: Data_out <= 16'h6BEE	;
				14'b01010111001001: Data_out <= 16'h6BE7	;
				14'b01010111001010: Data_out <= 16'h6BE0	;
				14'b01010111001011: Data_out <= 16'h6BD9	;
				14'b01010111001100: Data_out <= 16'h6BD2	;
				14'b01010111001101: Data_out <= 16'h6BCC	;
				14'b01010111001110: Data_out <= 16'h6BC5	;
				14'b01010111001111: Data_out <= 16'h6BBE	;
				14'b01010111010000: Data_out <= 16'h6BB7	;
				14'b01010111010001: Data_out <= 16'h6BB1	;
				14'b01010111010010: Data_out <= 16'h6BAA	;
				14'b01010111010011: Data_out <= 16'h6BA3	;
				14'b01010111010100: Data_out <= 16'h6B9C	;
				14'b01010111010101: Data_out <= 16'h6B95	;
				14'b01010111010110: Data_out <= 16'h6B8F	;
				14'b01010111010111: Data_out <= 16'h6B88	;
				14'b01010111011000: Data_out <= 16'h6B81	;
				14'b01010111011001: Data_out <= 16'h6B7A	;
				14'b01010111011010: Data_out <= 16'h6B73	;
				14'b01010111011011: Data_out <= 16'h6B6C	;
				14'b01010111011100: Data_out <= 16'h6B66	;
				14'b01010111011101: Data_out <= 16'h6B5F	;
				14'b01010111011110: Data_out <= 16'h6B58	;
				14'b01010111011111: Data_out <= 16'h6B51	;
				14'b01010111100000: Data_out <= 16'h6B4A	;
				14'b01010111100001: Data_out <= 16'h6B43	;
				14'b01010111100010: Data_out <= 16'h6B3C	;
				14'b01010111100011: Data_out <= 16'h6B36	;
				14'b01010111100100: Data_out <= 16'h6B2F	;
				14'b01010111100101: Data_out <= 16'h6B28	;
				14'b01010111100110: Data_out <= 16'h6B21	;
				14'b01010111100111: Data_out <= 16'h6B1A	;
				14'b01010111101000: Data_out <= 16'h6B13	;
				14'b01010111101001: Data_out <= 16'h6B0C	;
				14'b01010111101010: Data_out <= 16'h6B05	;
				14'b01010111101011: Data_out <= 16'h6AFF	;
				14'b01010111101100: Data_out <= 16'h6AF8	;
				14'b01010111101101: Data_out <= 16'h6AF1	;
				14'b01010111101110: Data_out <= 16'h6AEA	;
				14'b01010111101111: Data_out <= 16'h6AE3	;
				14'b01010111110000: Data_out <= 16'h6ADC	;
				14'b01010111110001: Data_out <= 16'h6AD5	;
				14'b01010111110010: Data_out <= 16'h6ACE	;
				14'b01010111110011: Data_out <= 16'h6AC7	;
				14'b01010111110100: Data_out <= 16'h6AC0	;
				14'b01010111110101: Data_out <= 16'h6AB9	;
				14'b01010111110110: Data_out <= 16'h6AB2	;
				14'b01010111110111: Data_out <= 16'h6AAC	;
				14'b01010111111000: Data_out <= 16'h6AA5	;
				14'b01010111111001: Data_out <= 16'h6A9E	;
				14'b01010111111010: Data_out <= 16'h6A97	;
				14'b01010111111011: Data_out <= 16'h6A90	;
				14'b01010111111100: Data_out <= 16'h6A89	;
				14'b01010111111101: Data_out <= 16'h6A82	;
				14'b01010111111110: Data_out <= 16'h6A7B	;
				14'b01010111111111: Data_out <= 16'h6A74	;
				14'b01011000000000: Data_out <= 16'h6A6D	;
				14'b01011000000001: Data_out <= 16'h6A66	;
				14'b01011000000010: Data_out <= 16'h6A5F	;
				14'b01011000000011: Data_out <= 16'h6A58	;
				14'b01011000000100: Data_out <= 16'h6A51	;
				14'b01011000000101: Data_out <= 16'h6A4A	;
				14'b01011000000110: Data_out <= 16'h6A43	;
				14'b01011000000111: Data_out <= 16'h6A3C	;
				14'b01011000001000: Data_out <= 16'h6A35	;
				14'b01011000001001: Data_out <= 16'h6A2E	;
				14'b01011000001010: Data_out <= 16'h6A27	;
				14'b01011000001011: Data_out <= 16'h6A20	;
				14'b01011000001100: Data_out <= 16'h6A19	;
				14'b01011000001101: Data_out <= 16'h6A12	;
				14'b01011000001110: Data_out <= 16'h6A0B	;
				14'b01011000001111: Data_out <= 16'h6A04	;
				14'b01011000010000: Data_out <= 16'h69FD	;
				14'b01011000010001: Data_out <= 16'h69F6	;
				14'b01011000010010: Data_out <= 16'h69EF	;
				14'b01011000010011: Data_out <= 16'h69E7	;
				14'b01011000010100: Data_out <= 16'h69E0	;
				14'b01011000010101: Data_out <= 16'h69D9	;
				14'b01011000010110: Data_out <= 16'h69D2	;
				14'b01011000010111: Data_out <= 16'h69CB	;
				14'b01011000011000: Data_out <= 16'h69C4	;
				14'b01011000011001: Data_out <= 16'h69BD	;
				14'b01011000011010: Data_out <= 16'h69B6	;
				14'b01011000011011: Data_out <= 16'h69AF	;
				14'b01011000011100: Data_out <= 16'h69A8	;
				14'b01011000011101: Data_out <= 16'h69A1	;
				14'b01011000011110: Data_out <= 16'h699A	;
				14'b01011000011111: Data_out <= 16'h6993	;
				14'b01011000100000: Data_out <= 16'h698B	;
				14'b01011000100001: Data_out <= 16'h6984	;
				14'b01011000100010: Data_out <= 16'h697D	;
				14'b01011000100011: Data_out <= 16'h6976	;
				14'b01011000100100: Data_out <= 16'h696F	;
				14'b01011000100101: Data_out <= 16'h6968	;
				14'b01011000100110: Data_out <= 16'h6961	;
				14'b01011000100111: Data_out <= 16'h695A	;
				14'b01011000101000: Data_out <= 16'h6952	;
				14'b01011000101001: Data_out <= 16'h694B	;
				14'b01011000101010: Data_out <= 16'h6944	;
				14'b01011000101011: Data_out <= 16'h693D	;
				14'b01011000101100: Data_out <= 16'h6936	;
				14'b01011000101101: Data_out <= 16'h692F	;
				14'b01011000101110: Data_out <= 16'h6928	;
				14'b01011000101111: Data_out <= 16'h6920	;
				14'b01011000110000: Data_out <= 16'h6919	;
				14'b01011000110001: Data_out <= 16'h6912	;
				14'b01011000110010: Data_out <= 16'h690B	;
				14'b01011000110011: Data_out <= 16'h6904	;
				14'b01011000110100: Data_out <= 16'h68FC	;
				14'b01011000110101: Data_out <= 16'h68F5	;
				14'b01011000110110: Data_out <= 16'h68EE	;
				14'b01011000110111: Data_out <= 16'h68E7	;
				14'b01011000111000: Data_out <= 16'h68E0	;
				14'b01011000111001: Data_out <= 16'h68D8	;
				14'b01011000111010: Data_out <= 16'h68D1	;
				14'b01011000111011: Data_out <= 16'h68CA	;
				14'b01011000111100: Data_out <= 16'h68C3	;
				14'b01011000111101: Data_out <= 16'h68BC	;
				14'b01011000111110: Data_out <= 16'h68B4	;
				14'b01011000111111: Data_out <= 16'h68AD	;
				14'b01011001000000: Data_out <= 16'h68A6	;
				14'b01011001000001: Data_out <= 16'h689F	;
				14'b01011001000010: Data_out <= 16'h6897	;
				14'b01011001000011: Data_out <= 16'h6890	;
				14'b01011001000100: Data_out <= 16'h6889	;
				14'b01011001000101: Data_out <= 16'h6882	;
				14'b01011001000110: Data_out <= 16'h687A	;
				14'b01011001000111: Data_out <= 16'h6873	;
				14'b01011001001000: Data_out <= 16'h686C	;
				14'b01011001001001: Data_out <= 16'h6865	;
				14'b01011001001010: Data_out <= 16'h685D	;
				14'b01011001001011: Data_out <= 16'h6856	;
				14'b01011001001100: Data_out <= 16'h684F	;
				14'b01011001001101: Data_out <= 16'h6848	;
				14'b01011001001110: Data_out <= 16'h6840	;
				14'b01011001001111: Data_out <= 16'h6839	;
				14'b01011001010000: Data_out <= 16'h6832	;
				14'b01011001010001: Data_out <= 16'h682A	;
				14'b01011001010010: Data_out <= 16'h6823	;
				14'b01011001010011: Data_out <= 16'h681C	;
				14'b01011001010100: Data_out <= 16'h6814	;
				14'b01011001010101: Data_out <= 16'h680D	;
				14'b01011001010110: Data_out <= 16'h6806	;
				14'b01011001010111: Data_out <= 16'h67FE	;
				14'b01011001011000: Data_out <= 16'h67F7	;
				14'b01011001011001: Data_out <= 16'h67F0	;
				14'b01011001011010: Data_out <= 16'h67E8	;
				14'b01011001011011: Data_out <= 16'h67E1	;
				14'b01011001011100: Data_out <= 16'h67DA	;
				14'b01011001011101: Data_out <= 16'h67D2	;
				14'b01011001011110: Data_out <= 16'h67CB	;
				14'b01011001011111: Data_out <= 16'h67C4	;
				14'b01011001100000: Data_out <= 16'h67BC	;
				14'b01011001100001: Data_out <= 16'h67B5	;
				14'b01011001100010: Data_out <= 16'h67AE	;
				14'b01011001100011: Data_out <= 16'h67A6	;
				14'b01011001100100: Data_out <= 16'h679F	;
				14'b01011001100101: Data_out <= 16'h6797	;
				14'b01011001100110: Data_out <= 16'h6790	;
				14'b01011001100111: Data_out <= 16'h6789	;
				14'b01011001101000: Data_out <= 16'h6781	;
				14'b01011001101001: Data_out <= 16'h677A	;
				14'b01011001101010: Data_out <= 16'h6773	;
				14'b01011001101011: Data_out <= 16'h676B	;
				14'b01011001101100: Data_out <= 16'h6764	;
				14'b01011001101101: Data_out <= 16'h675C	;
				14'b01011001101110: Data_out <= 16'h6755	;
				14'b01011001101111: Data_out <= 16'h674D	;
				14'b01011001110000: Data_out <= 16'h6746	;
				14'b01011001110001: Data_out <= 16'h673F	;
				14'b01011001110010: Data_out <= 16'h6737	;
				14'b01011001110011: Data_out <= 16'h6730	;
				14'b01011001110100: Data_out <= 16'h6728	;
				14'b01011001110101: Data_out <= 16'h6721	;
				14'b01011001110110: Data_out <= 16'h6719	;
				14'b01011001110111: Data_out <= 16'h6712	;
				14'b01011001111000: Data_out <= 16'h670B	;
				14'b01011001111001: Data_out <= 16'h6703	;
				14'b01011001111010: Data_out <= 16'h66FC	;
				14'b01011001111011: Data_out <= 16'h66F4	;
				14'b01011001111100: Data_out <= 16'h66ED	;
				14'b01011001111101: Data_out <= 16'h66E5	;
				14'b01011001111110: Data_out <= 16'h66DE	;
				14'b01011001111111: Data_out <= 16'h66D6	;
				14'b01011010000000: Data_out <= 16'h66CF	;
				14'b01011010000001: Data_out <= 16'h66C7	;
				14'b01011010000010: Data_out <= 16'h66C0	;
				14'b01011010000011: Data_out <= 16'h66B8	;
				14'b01011010000100: Data_out <= 16'h66B1	;
				14'b01011010000101: Data_out <= 16'h66A9	;
				14'b01011010000110: Data_out <= 16'h66A2	;
				14'b01011010000111: Data_out <= 16'h669A	;
				14'b01011010001000: Data_out <= 16'h6693	;
				14'b01011010001001: Data_out <= 16'h668B	;
				14'b01011010001010: Data_out <= 16'h6684	;
				14'b01011010001011: Data_out <= 16'h667C	;
				14'b01011010001100: Data_out <= 16'h6675	;
				14'b01011010001101: Data_out <= 16'h666D	;
				14'b01011010001110: Data_out <= 16'h6666	;
				14'b01011010001111: Data_out <= 16'h665E	;
				14'b01011010010000: Data_out <= 16'h6657	;
				14'b01011010010001: Data_out <= 16'h664F	;
				14'b01011010010010: Data_out <= 16'h6647	;
				14'b01011010010011: Data_out <= 16'h6640	;
				14'b01011010010100: Data_out <= 16'h6638	;
				14'b01011010010101: Data_out <= 16'h6631	;
				14'b01011010010110: Data_out <= 16'h6629	;
				14'b01011010010111: Data_out <= 16'h6622	;
				14'b01011010011000: Data_out <= 16'h661A	;
				14'b01011010011001: Data_out <= 16'h6612	;
				14'b01011010011010: Data_out <= 16'h660B	;
				14'b01011010011011: Data_out <= 16'h6603	;
				14'b01011010011100: Data_out <= 16'h65FC	;
				14'b01011010011101: Data_out <= 16'h65F4	;
				14'b01011010011110: Data_out <= 16'h65EC	;
				14'b01011010011111: Data_out <= 16'h65E5	;
				14'b01011010100000: Data_out <= 16'h65DD	;
				14'b01011010100001: Data_out <= 16'h65D6	;
				14'b01011010100010: Data_out <= 16'h65CE	;
				14'b01011010100011: Data_out <= 16'h65C6	;
				14'b01011010100100: Data_out <= 16'h65BF	;
				14'b01011010100101: Data_out <= 16'h65B7	;
				14'b01011010100110: Data_out <= 16'h65B0	;
				14'b01011010100111: Data_out <= 16'h65A8	;
				14'b01011010101000: Data_out <= 16'h65A0	;
				14'b01011010101001: Data_out <= 16'h6599	;
				14'b01011010101010: Data_out <= 16'h6591	;
				14'b01011010101011: Data_out <= 16'h6589	;
				14'b01011010101100: Data_out <= 16'h6582	;
				14'b01011010101101: Data_out <= 16'h657A	;
				14'b01011010101110: Data_out <= 16'h6572	;
				14'b01011010101111: Data_out <= 16'h656B	;
				14'b01011010110000: Data_out <= 16'h6563	;
				14'b01011010110001: Data_out <= 16'h655B	;
				14'b01011010110010: Data_out <= 16'h6554	;
				14'b01011010110011: Data_out <= 16'h654C	;
				14'b01011010110100: Data_out <= 16'h6544	;
				14'b01011010110101: Data_out <= 16'h653D	;
				14'b01011010110110: Data_out <= 16'h6535	;
				14'b01011010110111: Data_out <= 16'h652D	;
				14'b01011010111000: Data_out <= 16'h6526	;
				14'b01011010111001: Data_out <= 16'h651E	;
				14'b01011010111010: Data_out <= 16'h6516	;
				14'b01011010111011: Data_out <= 16'h650E	;
				14'b01011010111100: Data_out <= 16'h6507	;
				14'b01011010111101: Data_out <= 16'h64FF	;
				14'b01011010111110: Data_out <= 16'h64F7	;
				14'b01011010111111: Data_out <= 16'h64F0	;
				14'b01011011000000: Data_out <= 16'h64E8	;
				14'b01011011000001: Data_out <= 16'h64E0	;
				14'b01011011000010: Data_out <= 16'h64D8	;
				14'b01011011000011: Data_out <= 16'h64D1	;
				14'b01011011000100: Data_out <= 16'h64C9	;
				14'b01011011000101: Data_out <= 16'h64C1	;
				14'b01011011000110: Data_out <= 16'h64B9	;
				14'b01011011000111: Data_out <= 16'h64B2	;
				14'b01011011001000: Data_out <= 16'h64AA	;
				14'b01011011001001: Data_out <= 16'h64A2	;
				14'b01011011001010: Data_out <= 16'h649A	;
				14'b01011011001011: Data_out <= 16'h6493	;
				14'b01011011001100: Data_out <= 16'h648B	;
				14'b01011011001101: Data_out <= 16'h6483	;
				14'b01011011001110: Data_out <= 16'h647B	;
				14'b01011011001111: Data_out <= 16'h6473	;
				14'b01011011010000: Data_out <= 16'h646C	;
				14'b01011011010001: Data_out <= 16'h6464	;
				14'b01011011010010: Data_out <= 16'h645C	;
				14'b01011011010011: Data_out <= 16'h6454	;
				14'b01011011010100: Data_out <= 16'h644C	;
				14'b01011011010101: Data_out <= 16'h6445	;
				14'b01011011010110: Data_out <= 16'h643D	;
				14'b01011011010111: Data_out <= 16'h6435	;
				14'b01011011011000: Data_out <= 16'h642D	;
				14'b01011011011001: Data_out <= 16'h6425	;
				14'b01011011011010: Data_out <= 16'h641E	;
				14'b01011011011011: Data_out <= 16'h6416	;
				14'b01011011011100: Data_out <= 16'h640E	;
				14'b01011011011101: Data_out <= 16'h6406	;
				14'b01011011011110: Data_out <= 16'h63FE	;
				14'b01011011011111: Data_out <= 16'h63F6	;
				14'b01011011100000: Data_out <= 16'h63EF	;
				14'b01011011100001: Data_out <= 16'h63E7	;
				14'b01011011100010: Data_out <= 16'h63DF	;
				14'b01011011100011: Data_out <= 16'h63D7	;
				14'b01011011100100: Data_out <= 16'h63CF	;
				14'b01011011100101: Data_out <= 16'h63C7	;
				14'b01011011100110: Data_out <= 16'h63BF	;
				14'b01011011100111: Data_out <= 16'h63B7	;
				14'b01011011101000: Data_out <= 16'h63B0	;
				14'b01011011101001: Data_out <= 16'h63A8	;
				14'b01011011101010: Data_out <= 16'h63A0	;
				14'b01011011101011: Data_out <= 16'h6398	;
				14'b01011011101100: Data_out <= 16'h6390	;
				14'b01011011101101: Data_out <= 16'h6388	;
				14'b01011011101110: Data_out <= 16'h6380	;
				14'b01011011101111: Data_out <= 16'h6378	;
				14'b01011011110000: Data_out <= 16'h6370	;
				14'b01011011110001: Data_out <= 16'h6368	;
				14'b01011011110010: Data_out <= 16'h6361	;
				14'b01011011110011: Data_out <= 16'h6359	;
				14'b01011011110100: Data_out <= 16'h6351	;
				14'b01011011110101: Data_out <= 16'h6349	;
				14'b01011011110110: Data_out <= 16'h6341	;
				14'b01011011110111: Data_out <= 16'h6339	;
				14'b01011011111000: Data_out <= 16'h6331	;
				14'b01011011111001: Data_out <= 16'h6329	;
				14'b01011011111010: Data_out <= 16'h6321	;
				14'b01011011111011: Data_out <= 16'h6319	;
				14'b01011011111100: Data_out <= 16'h6311	;
				14'b01011011111101: Data_out <= 16'h6309	;
				14'b01011011111110: Data_out <= 16'h6301	;
				14'b01011011111111: Data_out <= 16'h62F9	;
				14'b01011100000000: Data_out <= 16'h62F1	;
				14'b01011100000001: Data_out <= 16'h62E9	;
				14'b01011100000010: Data_out <= 16'h62E1	;
				14'b01011100000011: Data_out <= 16'h62D9	;
				14'b01011100000100: Data_out <= 16'h62D1	;
				14'b01011100000101: Data_out <= 16'h62C9	;
				14'b01011100000110: Data_out <= 16'h62C1	;
				14'b01011100000111: Data_out <= 16'h62B9	;
				14'b01011100001000: Data_out <= 16'h62B1	;
				14'b01011100001001: Data_out <= 16'h62A9	;
				14'b01011100001010: Data_out <= 16'h62A1	;
				14'b01011100001011: Data_out <= 16'h6299	;
				14'b01011100001100: Data_out <= 16'h6291	;
				14'b01011100001101: Data_out <= 16'h6289	;
				14'b01011100001110: Data_out <= 16'h6281	;
				14'b01011100001111: Data_out <= 16'h6279	;
				14'b01011100010000: Data_out <= 16'h6271	;
				14'b01011100010001: Data_out <= 16'h6269	;
				14'b01011100010010: Data_out <= 16'h6261	;
				14'b01011100010011: Data_out <= 16'h6259	;
				14'b01011100010100: Data_out <= 16'h6251	;
				14'b01011100010101: Data_out <= 16'h6249	;
				14'b01011100010110: Data_out <= 16'h6241	;
				14'b01011100010111: Data_out <= 16'h6239	;
				14'b01011100011000: Data_out <= 16'h6231	;
				14'b01011100011001: Data_out <= 16'h6229	;
				14'b01011100011010: Data_out <= 16'h6221	;
				14'b01011100011011: Data_out <= 16'h6219	;
				14'b01011100011100: Data_out <= 16'h6211	;
				14'b01011100011101: Data_out <= 16'h6209	;
				14'b01011100011110: Data_out <= 16'h6201	;
				14'b01011100011111: Data_out <= 16'h61F8	;
				14'b01011100100000: Data_out <= 16'h61F0	;
				14'b01011100100001: Data_out <= 16'h61E8	;
				14'b01011100100010: Data_out <= 16'h61E0	;
				14'b01011100100011: Data_out <= 16'h61D8	;
				14'b01011100100100: Data_out <= 16'h61D0	;
				14'b01011100100101: Data_out <= 16'h61C8	;
				14'b01011100100110: Data_out <= 16'h61C0	;
				14'b01011100100111: Data_out <= 16'h61B8	;
				14'b01011100101000: Data_out <= 16'h61AF	;
				14'b01011100101001: Data_out <= 16'h61A7	;
				14'b01011100101010: Data_out <= 16'h619F	;
				14'b01011100101011: Data_out <= 16'h6197	;
				14'b01011100101100: Data_out <= 16'h618F	;
				14'b01011100101101: Data_out <= 16'h6187	;
				14'b01011100101110: Data_out <= 16'h617F	;
				14'b01011100101111: Data_out <= 16'h6177	;
				14'b01011100110000: Data_out <= 16'h616E	;
				14'b01011100110001: Data_out <= 16'h6166	;
				14'b01011100110010: Data_out <= 16'h615E	;
				14'b01011100110011: Data_out <= 16'h6156	;
				14'b01011100110100: Data_out <= 16'h614E	;
				14'b01011100110101: Data_out <= 16'h6146	;
				14'b01011100110110: Data_out <= 16'h613D	;
				14'b01011100110111: Data_out <= 16'h6135	;
				14'b01011100111000: Data_out <= 16'h612D	;
				14'b01011100111001: Data_out <= 16'h6125	;
				14'b01011100111010: Data_out <= 16'h611D	;
				14'b01011100111011: Data_out <= 16'h6115	;
				14'b01011100111100: Data_out <= 16'h610C	;
				14'b01011100111101: Data_out <= 16'h6104	;
				14'b01011100111110: Data_out <= 16'h60FC	;
				14'b01011100111111: Data_out <= 16'h60F4	;
				14'b01011101000000: Data_out <= 16'h60EC	;
				14'b01011101000001: Data_out <= 16'h60E3	;
				14'b01011101000010: Data_out <= 16'h60DB	;
				14'b01011101000011: Data_out <= 16'h60D3	;
				14'b01011101000100: Data_out <= 16'h60CB	;
				14'b01011101000101: Data_out <= 16'h60C2	;
				14'b01011101000110: Data_out <= 16'h60BA	;
				14'b01011101000111: Data_out <= 16'h60B2	;
				14'b01011101001000: Data_out <= 16'h60AA	;
				14'b01011101001001: Data_out <= 16'h60A2	;
				14'b01011101001010: Data_out <= 16'h6099	;
				14'b01011101001011: Data_out <= 16'h6091	;
				14'b01011101001100: Data_out <= 16'h6089	;
				14'b01011101001101: Data_out <= 16'h6081	;
				14'b01011101001110: Data_out <= 16'h6078	;
				14'b01011101001111: Data_out <= 16'h6070	;
				14'b01011101010000: Data_out <= 16'h6068	;
				14'b01011101010001: Data_out <= 16'h6060	;
				14'b01011101010010: Data_out <= 16'h6057	;
				14'b01011101010011: Data_out <= 16'h604F	;
				14'b01011101010100: Data_out <= 16'h6047	;
				14'b01011101010101: Data_out <= 16'h603E	;
				14'b01011101010110: Data_out <= 16'h6036	;
				14'b01011101010111: Data_out <= 16'h602E	;
				14'b01011101011000: Data_out <= 16'h6026	;
				14'b01011101011001: Data_out <= 16'h601D	;
				14'b01011101011010: Data_out <= 16'h6015	;
				14'b01011101011011: Data_out <= 16'h600D	;
				14'b01011101011100: Data_out <= 16'h6004	;
				14'b01011101011101: Data_out <= 16'h5FFC	;
				14'b01011101011110: Data_out <= 16'h5FF4	;
				14'b01011101011111: Data_out <= 16'h5FEB	;
				14'b01011101100000: Data_out <= 16'h5FE3	;
				14'b01011101100001: Data_out <= 16'h5FDB	;
				14'b01011101100010: Data_out <= 16'h5FD2	;
				14'b01011101100011: Data_out <= 16'h5FCA	;
				14'b01011101100100: Data_out <= 16'h5FC2	;
				14'b01011101100101: Data_out <= 16'h5FB9	;
				14'b01011101100110: Data_out <= 16'h5FB1	;
				14'b01011101100111: Data_out <= 16'h5FA9	;
				14'b01011101101000: Data_out <= 16'h5FA0	;
				14'b01011101101001: Data_out <= 16'h5F98	;
				14'b01011101101010: Data_out <= 16'h5F90	;
				14'b01011101101011: Data_out <= 16'h5F87	;
				14'b01011101101100: Data_out <= 16'h5F7F	;
				14'b01011101101101: Data_out <= 16'h5F77	;
				14'b01011101101110: Data_out <= 16'h5F6E	;
				14'b01011101101111: Data_out <= 16'h5F66	;
				14'b01011101110000: Data_out <= 16'h5F5D	;
				14'b01011101110001: Data_out <= 16'h5F55	;
				14'b01011101110010: Data_out <= 16'h5F4D	;
				14'b01011101110011: Data_out <= 16'h5F44	;
				14'b01011101110100: Data_out <= 16'h5F3C	;
				14'b01011101110101: Data_out <= 16'h5F33	;
				14'b01011101110110: Data_out <= 16'h5F2B	;
				14'b01011101110111: Data_out <= 16'h5F23	;
				14'b01011101111000: Data_out <= 16'h5F1A	;
				14'b01011101111001: Data_out <= 16'h5F12	;
				14'b01011101111010: Data_out <= 16'h5F09	;
				14'b01011101111011: Data_out <= 16'h5F01	;
				14'b01011101111100: Data_out <= 16'h5EF9	;
				14'b01011101111101: Data_out <= 16'h5EF0	;
				14'b01011101111110: Data_out <= 16'h5EE8	;
				14'b01011101111111: Data_out <= 16'h5EDF	;
				14'b01011110000000: Data_out <= 16'h5ED7	;
				14'b01011110000001: Data_out <= 16'h5ECE	;
				14'b01011110000010: Data_out <= 16'h5EC6	;
				14'b01011110000011: Data_out <= 16'h5EBE	;
				14'b01011110000100: Data_out <= 16'h5EB5	;
				14'b01011110000101: Data_out <= 16'h5EAD	;
				14'b01011110000110: Data_out <= 16'h5EA4	;
				14'b01011110000111: Data_out <= 16'h5E9C	;
				14'b01011110001000: Data_out <= 16'h5E93	;
				14'b01011110001001: Data_out <= 16'h5E8B	;
				14'b01011110001010: Data_out <= 16'h5E82	;
				14'b01011110001011: Data_out <= 16'h5E7A	;
				14'b01011110001100: Data_out <= 16'h5E71	;
				14'b01011110001101: Data_out <= 16'h5E69	;
				14'b01011110001110: Data_out <= 16'h5E60	;
				14'b01011110001111: Data_out <= 16'h5E58	;
				14'b01011110010000: Data_out <= 16'h5E4F	;
				14'b01011110010001: Data_out <= 16'h5E47	;
				14'b01011110010010: Data_out <= 16'h5E3E	;
				14'b01011110010011: Data_out <= 16'h5E36	;
				14'b01011110010100: Data_out <= 16'h5E2D	;
				14'b01011110010101: Data_out <= 16'h5E25	;
				14'b01011110010110: Data_out <= 16'h5E1C	;
				14'b01011110010111: Data_out <= 16'h5E14	;
				14'b01011110011000: Data_out <= 16'h5E0B	;
				14'b01011110011001: Data_out <= 16'h5E03	;
				14'b01011110011010: Data_out <= 16'h5DFA	;
				14'b01011110011011: Data_out <= 16'h5DF2	;
				14'b01011110011100: Data_out <= 16'h5DE9	;
				14'b01011110011101: Data_out <= 16'h5DE1	;
				14'b01011110011110: Data_out <= 16'h5DD8	;
				14'b01011110011111: Data_out <= 16'h5DD0	;
				14'b01011110100000: Data_out <= 16'h5DC7	;
				14'b01011110100001: Data_out <= 16'h5DBE	;
				14'b01011110100010: Data_out <= 16'h5DB6	;
				14'b01011110100011: Data_out <= 16'h5DAD	;
				14'b01011110100100: Data_out <= 16'h5DA5	;
				14'b01011110100101: Data_out <= 16'h5D9C	;
				14'b01011110100110: Data_out <= 16'h5D94	;
				14'b01011110100111: Data_out <= 16'h5D8B	;
				14'b01011110101000: Data_out <= 16'h5D82	;
				14'b01011110101001: Data_out <= 16'h5D7A	;
				14'b01011110101010: Data_out <= 16'h5D71	;
				14'b01011110101011: Data_out <= 16'h5D69	;
				14'b01011110101100: Data_out <= 16'h5D60	;
				14'b01011110101101: Data_out <= 16'h5D58	;
				14'b01011110101110: Data_out <= 16'h5D4F	;
				14'b01011110101111: Data_out <= 16'h5D46	;
				14'b01011110110000: Data_out <= 16'h5D3E	;
				14'b01011110110001: Data_out <= 16'h5D35	;
				14'b01011110110010: Data_out <= 16'h5D2C	;
				14'b01011110110011: Data_out <= 16'h5D24	;
				14'b01011110110100: Data_out <= 16'h5D1B	;
				14'b01011110110101: Data_out <= 16'h5D13	;
				14'b01011110110110: Data_out <= 16'h5D0A	;
				14'b01011110110111: Data_out <= 16'h5D01	;
				14'b01011110111000: Data_out <= 16'h5CF9	;
				14'b01011110111001: Data_out <= 16'h5CF0	;
				14'b01011110111010: Data_out <= 16'h5CE7	;
				14'b01011110111011: Data_out <= 16'h5CDF	;
				14'b01011110111100: Data_out <= 16'h5CD6	;
				14'b01011110111101: Data_out <= 16'h5CCD	;
				14'b01011110111110: Data_out <= 16'h5CC5	;
				14'b01011110111111: Data_out <= 16'h5CBC	;
				14'b01011111000000: Data_out <= 16'h5CB4	;
				14'b01011111000001: Data_out <= 16'h5CAB	;
				14'b01011111000010: Data_out <= 16'h5CA2	;
				14'b01011111000011: Data_out <= 16'h5C99	;
				14'b01011111000100: Data_out <= 16'h5C91	;
				14'b01011111000101: Data_out <= 16'h5C88	;
				14'b01011111000110: Data_out <= 16'h5C7F	;
				14'b01011111000111: Data_out <= 16'h5C77	;
				14'b01011111001000: Data_out <= 16'h5C6E	;
				14'b01011111001001: Data_out <= 16'h5C65	;
				14'b01011111001010: Data_out <= 16'h5C5D	;
				14'b01011111001011: Data_out <= 16'h5C54	;
				14'b01011111001100: Data_out <= 16'h5C4B	;
				14'b01011111001101: Data_out <= 16'h5C43	;
				14'b01011111001110: Data_out <= 16'h5C3A	;
				14'b01011111001111: Data_out <= 16'h5C31	;
				14'b01011111010000: Data_out <= 16'h5C28	;
				14'b01011111010001: Data_out <= 16'h5C20	;
				14'b01011111010010: Data_out <= 16'h5C17	;
				14'b01011111010011: Data_out <= 16'h5C0E	;
				14'b01011111010100: Data_out <= 16'h5C06	;
				14'b01011111010101: Data_out <= 16'h5BFD	;
				14'b01011111010110: Data_out <= 16'h5BF4	;
				14'b01011111010111: Data_out <= 16'h5BEB	;
				14'b01011111011000: Data_out <= 16'h5BE3	;
				14'b01011111011001: Data_out <= 16'h5BDA	;
				14'b01011111011010: Data_out <= 16'h5BD1	;
				14'b01011111011011: Data_out <= 16'h5BC8	;
				14'b01011111011100: Data_out <= 16'h5BC0	;
				14'b01011111011101: Data_out <= 16'h5BB7	;
				14'b01011111011110: Data_out <= 16'h5BAE	;
				14'b01011111011111: Data_out <= 16'h5BA5	;
				14'b01011111100000: Data_out <= 16'h5B9C	;
				14'b01011111100001: Data_out <= 16'h5B94	;
				14'b01011111100010: Data_out <= 16'h5B8B	;
				14'b01011111100011: Data_out <= 16'h5B82	;
				14'b01011111100100: Data_out <= 16'h5B79	;
				14'b01011111100101: Data_out <= 16'h5B71	;
				14'b01011111100110: Data_out <= 16'h5B68	;
				14'b01011111100111: Data_out <= 16'h5B5F	;
				14'b01011111101000: Data_out <= 16'h5B56	;
				14'b01011111101001: Data_out <= 16'h5B4D	;
				14'b01011111101010: Data_out <= 16'h5B45	;
				14'b01011111101011: Data_out <= 16'h5B3C	;
				14'b01011111101100: Data_out <= 16'h5B33	;
				14'b01011111101101: Data_out <= 16'h5B2A	;
				14'b01011111101110: Data_out <= 16'h5B21	;
				14'b01011111101111: Data_out <= 16'h5B18	;
				14'b01011111110000: Data_out <= 16'h5B10	;
				14'b01011111110001: Data_out <= 16'h5B07	;
				14'b01011111110010: Data_out <= 16'h5AFE	;
				14'b01011111110011: Data_out <= 16'h5AF5	;
				14'b01011111110100: Data_out <= 16'h5AEC	;
				14'b01011111110101: Data_out <= 16'h5AE3	;
				14'b01011111110110: Data_out <= 16'h5ADB	;
				14'b01011111110111: Data_out <= 16'h5AD2	;
				14'b01011111111000: Data_out <= 16'h5AC9	;
				14'b01011111111001: Data_out <= 16'h5AC0	;
				14'b01011111111010: Data_out <= 16'h5AB7	;
				14'b01011111111011: Data_out <= 16'h5AAE	;
				14'b01011111111100: Data_out <= 16'h5AA5	;
				14'b01011111111101: Data_out <= 16'h5A9D	;
				14'b01011111111110: Data_out <= 16'h5A94	;
				14'b01011111111111: Data_out <= 16'h5A8B	;
				14'b01100000000000: Data_out <= 16'h5A82	;
				14'b01100000000001: Data_out <= 16'h5A79	;
				14'b01100000000010: Data_out <= 16'h5A70	;
				14'b01100000000011: Data_out <= 16'h5A67	;
				14'b01100000000100: Data_out <= 16'h5A5E	;
				14'b01100000000101: Data_out <= 16'h5A55	;
				14'b01100000000110: Data_out <= 16'h5A4C	;
				14'b01100000000111: Data_out <= 16'h5A44	;
				14'b01100000001000: Data_out <= 16'h5A3B	;
				14'b01100000001001: Data_out <= 16'h5A32	;
				14'b01100000001010: Data_out <= 16'h5A29	;
				14'b01100000001011: Data_out <= 16'h5A20	;
				14'b01100000001100: Data_out <= 16'h5A17	;
				14'b01100000001101: Data_out <= 16'h5A0E	;
				14'b01100000001110: Data_out <= 16'h5A05	;
				14'b01100000001111: Data_out <= 16'h59FC	;
				14'b01100000010000: Data_out <= 16'h59F3	;
				14'b01100000010001: Data_out <= 16'h59EA	;
				14'b01100000010010: Data_out <= 16'h59E1	;
				14'b01100000010011: Data_out <= 16'h59D8	;
				14'b01100000010100: Data_out <= 16'h59CF	;
				14'b01100000010101: Data_out <= 16'h59C7	;
				14'b01100000010110: Data_out <= 16'h59BE	;
				14'b01100000010111: Data_out <= 16'h59B5	;
				14'b01100000011000: Data_out <= 16'h59AC	;
				14'b01100000011001: Data_out <= 16'h59A3	;
				14'b01100000011010: Data_out <= 16'h599A	;
				14'b01100000011011: Data_out <= 16'h5991	;
				14'b01100000011100: Data_out <= 16'h5988	;
				14'b01100000011101: Data_out <= 16'h597F	;
				14'b01100000011110: Data_out <= 16'h5976	;
				14'b01100000011111: Data_out <= 16'h596D	;
				14'b01100000100000: Data_out <= 16'h5964	;
				14'b01100000100001: Data_out <= 16'h595B	;
				14'b01100000100010: Data_out <= 16'h5952	;
				14'b01100000100011: Data_out <= 16'h5949	;
				14'b01100000100100: Data_out <= 16'h5940	;
				14'b01100000100101: Data_out <= 16'h5937	;
				14'b01100000100110: Data_out <= 16'h592E	;
				14'b01100000100111: Data_out <= 16'h5925	;
				14'b01100000101000: Data_out <= 16'h591C	;
				14'b01100000101001: Data_out <= 16'h5913	;
				14'b01100000101010: Data_out <= 16'h590A	;
				14'b01100000101011: Data_out <= 16'h5901	;
				14'b01100000101100: Data_out <= 16'h58F8	;
				14'b01100000101101: Data_out <= 16'h58EF	;
				14'b01100000101110: Data_out <= 16'h58E6	;
				14'b01100000101111: Data_out <= 16'h58DD	;
				14'b01100000110000: Data_out <= 16'h58D3	;
				14'b01100000110001: Data_out <= 16'h58CA	;
				14'b01100000110010: Data_out <= 16'h58C1	;
				14'b01100000110011: Data_out <= 16'h58B8	;
				14'b01100000110100: Data_out <= 16'h58AF	;
				14'b01100000110101: Data_out <= 16'h58A6	;
				14'b01100000110110: Data_out <= 16'h589D	;
				14'b01100000110111: Data_out <= 16'h5894	;
				14'b01100000111000: Data_out <= 16'h588B	;
				14'b01100000111001: Data_out <= 16'h5882	;
				14'b01100000111010: Data_out <= 16'h5879	;
				14'b01100000111011: Data_out <= 16'h5870	;
				14'b01100000111100: Data_out <= 16'h5867	;
				14'b01100000111101: Data_out <= 16'h585E	;
				14'b01100000111110: Data_out <= 16'h5854	;
				14'b01100000111111: Data_out <= 16'h584B	;
				14'b01100001000000: Data_out <= 16'h5842	;
				14'b01100001000001: Data_out <= 16'h5839	;
				14'b01100001000010: Data_out <= 16'h5830	;
				14'b01100001000011: Data_out <= 16'h5827	;
				14'b01100001000100: Data_out <= 16'h581E	;
				14'b01100001000101: Data_out <= 16'h5815	;
				14'b01100001000110: Data_out <= 16'h580C	;
				14'b01100001000111: Data_out <= 16'h5802	;
				14'b01100001001000: Data_out <= 16'h57F9	;
				14'b01100001001001: Data_out <= 16'h57F0	;
				14'b01100001001010: Data_out <= 16'h57E7	;
				14'b01100001001011: Data_out <= 16'h57DE	;
				14'b01100001001100: Data_out <= 16'h57D5	;
				14'b01100001001101: Data_out <= 16'h57CC	;
				14'b01100001001110: Data_out <= 16'h57C3	;
				14'b01100001001111: Data_out <= 16'h57B9	;
				14'b01100001010000: Data_out <= 16'h57B0	;
				14'b01100001010001: Data_out <= 16'h57A7	;
				14'b01100001010010: Data_out <= 16'h579E	;
				14'b01100001010011: Data_out <= 16'h5795	;
				14'b01100001010100: Data_out <= 16'h578C	;
				14'b01100001010101: Data_out <= 16'h5782	;
				14'b01100001010110: Data_out <= 16'h5779	;
				14'b01100001010111: Data_out <= 16'h5770	;
				14'b01100001011000: Data_out <= 16'h5767	;
				14'b01100001011001: Data_out <= 16'h575E	;
				14'b01100001011010: Data_out <= 16'h5755	;
				14'b01100001011011: Data_out <= 16'h574B	;
				14'b01100001011100: Data_out <= 16'h5742	;
				14'b01100001011101: Data_out <= 16'h5739	;
				14'b01100001011110: Data_out <= 16'h5730	;
				14'b01100001011111: Data_out <= 16'h5727	;
				14'b01100001100000: Data_out <= 16'h571D	;
				14'b01100001100001: Data_out <= 16'h5714	;
				14'b01100001100010: Data_out <= 16'h570B	;
				14'b01100001100011: Data_out <= 16'h5702	;
				14'b01100001100100: Data_out <= 16'h56F9	;
				14'b01100001100101: Data_out <= 16'h56EF	;
				14'b01100001100110: Data_out <= 16'h56E6	;
				14'b01100001100111: Data_out <= 16'h56DD	;
				14'b01100001101000: Data_out <= 16'h56D4	;
				14'b01100001101001: Data_out <= 16'h56CA	;
				14'b01100001101010: Data_out <= 16'h56C1	;
				14'b01100001101011: Data_out <= 16'h56B8	;
				14'b01100001101100: Data_out <= 16'h56AF	;
				14'b01100001101101: Data_out <= 16'h56A5	;
				14'b01100001101110: Data_out <= 16'h569C	;
				14'b01100001101111: Data_out <= 16'h5693	;
				14'b01100001110000: Data_out <= 16'h568A	;
				14'b01100001110001: Data_out <= 16'h5680	;
				14'b01100001110010: Data_out <= 16'h5677	;
				14'b01100001110011: Data_out <= 16'h566E	;
				14'b01100001110100: Data_out <= 16'h5665	;
				14'b01100001110101: Data_out <= 16'h565B	;
				14'b01100001110110: Data_out <= 16'h5652	;
				14'b01100001110111: Data_out <= 16'h5649	;
				14'b01100001111000: Data_out <= 16'h563F	;
				14'b01100001111001: Data_out <= 16'h5636	;
				14'b01100001111010: Data_out <= 16'h562D	;
				14'b01100001111011: Data_out <= 16'h5624	;
				14'b01100001111100: Data_out <= 16'h561A	;
				14'b01100001111101: Data_out <= 16'h5611	;
				14'b01100001111110: Data_out <= 16'h5608	;
				14'b01100001111111: Data_out <= 16'h55FE	;
				14'b01100010000000: Data_out <= 16'h55F5	;
				14'b01100010000001: Data_out <= 16'h55EC	;
				14'b01100010000010: Data_out <= 16'h55E2	;
				14'b01100010000011: Data_out <= 16'h55D9	;
				14'b01100010000100: Data_out <= 16'h55D0	;
				14'b01100010000101: Data_out <= 16'h55C6	;
				14'b01100010000110: Data_out <= 16'h55BD	;
				14'b01100010000111: Data_out <= 16'h55B4	;
				14'b01100010001000: Data_out <= 16'h55AA	;
				14'b01100010001001: Data_out <= 16'h55A1	;
				14'b01100010001010: Data_out <= 16'h5598	;
				14'b01100010001011: Data_out <= 16'h558E	;
				14'b01100010001100: Data_out <= 16'h5585	;
				14'b01100010001101: Data_out <= 16'h557C	;
				14'b01100010001110: Data_out <= 16'h5572	;
				14'b01100010001111: Data_out <= 16'h5569	;
				14'b01100010010000: Data_out <= 16'h5560	;
				14'b01100010010001: Data_out <= 16'h5556	;
				14'b01100010010010: Data_out <= 16'h554D	;
				14'b01100010010011: Data_out <= 16'h5544	;
				14'b01100010010100: Data_out <= 16'h553A	;
				14'b01100010010101: Data_out <= 16'h5531	;
				14'b01100010010110: Data_out <= 16'h5527	;
				14'b01100010010111: Data_out <= 16'h551E	;
				14'b01100010011000: Data_out <= 16'h5515	;
				14'b01100010011001: Data_out <= 16'h550B	;
				14'b01100010011010: Data_out <= 16'h5502	;
				14'b01100010011011: Data_out <= 16'h54F9	;
				14'b01100010011100: Data_out <= 16'h54EF	;
				14'b01100010011101: Data_out <= 16'h54E6	;
				14'b01100010011110: Data_out <= 16'h54DC	;
				14'b01100010011111: Data_out <= 16'h54D3	;
				14'b01100010100000: Data_out <= 16'h54C9	;
				14'b01100010100001: Data_out <= 16'h54C0	;
				14'b01100010100010: Data_out <= 16'h54B7	;
				14'b01100010100011: Data_out <= 16'h54AD	;
				14'b01100010100100: Data_out <= 16'h54A4	;
				14'b01100010100101: Data_out <= 16'h549A	;
				14'b01100010100110: Data_out <= 16'h5491	;
				14'b01100010100111: Data_out <= 16'h5488	;
				14'b01100010101000: Data_out <= 16'h547E	;
				14'b01100010101001: Data_out <= 16'h5475	;
				14'b01100010101010: Data_out <= 16'h546B	;
				14'b01100010101011: Data_out <= 16'h5462	;
				14'b01100010101100: Data_out <= 16'h5458	;
				14'b01100010101101: Data_out <= 16'h544F	;
				14'b01100010101110: Data_out <= 16'h5445	;
				14'b01100010101111: Data_out <= 16'h543C	;
				14'b01100010110000: Data_out <= 16'h5432	;
				14'b01100010110001: Data_out <= 16'h5429	;
				14'b01100010110010: Data_out <= 16'h5420	;
				14'b01100010110011: Data_out <= 16'h5416	;
				14'b01100010110100: Data_out <= 16'h540D	;
				14'b01100010110101: Data_out <= 16'h5403	;
				14'b01100010110110: Data_out <= 16'h53FA	;
				14'b01100010110111: Data_out <= 16'h53F0	;
				14'b01100010111000: Data_out <= 16'h53E7	;
				14'b01100010111001: Data_out <= 16'h53DD	;
				14'b01100010111010: Data_out <= 16'h53D4	;
				14'b01100010111011: Data_out <= 16'h53CA	;
				14'b01100010111100: Data_out <= 16'h53C1	;
				14'b01100010111101: Data_out <= 16'h53B7	;
				14'b01100010111110: Data_out <= 16'h53AE	;
				14'b01100010111111: Data_out <= 16'h53A4	;
				14'b01100011000000: Data_out <= 16'h539B	;
				14'b01100011000001: Data_out <= 16'h5391	;
				14'b01100011000010: Data_out <= 16'h5388	;
				14'b01100011000011: Data_out <= 16'h537E	;
				14'b01100011000100: Data_out <= 16'h5375	;
				14'b01100011000101: Data_out <= 16'h536B	;
				14'b01100011000110: Data_out <= 16'h5361	;
				14'b01100011000111: Data_out <= 16'h5358	;
				14'b01100011001000: Data_out <= 16'h534E	;
				14'b01100011001001: Data_out <= 16'h5345	;
				14'b01100011001010: Data_out <= 16'h533B	;
				14'b01100011001011: Data_out <= 16'h5332	;
				14'b01100011001100: Data_out <= 16'h5328	;
				14'b01100011001101: Data_out <= 16'h531F	;
				14'b01100011001110: Data_out <= 16'h5315	;
				14'b01100011001111: Data_out <= 16'h530C	;
				14'b01100011010000: Data_out <= 16'h5302	;
				14'b01100011010001: Data_out <= 16'h52F8	;
				14'b01100011010010: Data_out <= 16'h52EF	;
				14'b01100011010011: Data_out <= 16'h52E5	;
				14'b01100011010100: Data_out <= 16'h52DC	;
				14'b01100011010101: Data_out <= 16'h52D2	;
				14'b01100011010110: Data_out <= 16'h52C9	;
				14'b01100011010111: Data_out <= 16'h52BF	;
				14'b01100011011000: Data_out <= 16'h52B5	;
				14'b01100011011001: Data_out <= 16'h52AC	;
				14'b01100011011010: Data_out <= 16'h52A2	;
				14'b01100011011011: Data_out <= 16'h5299	;
				14'b01100011011100: Data_out <= 16'h528F	;
				14'b01100011011101: Data_out <= 16'h5285	;
				14'b01100011011110: Data_out <= 16'h527C	;
				14'b01100011011111: Data_out <= 16'h5272	;
				14'b01100011100000: Data_out <= 16'h5269	;
				14'b01100011100001: Data_out <= 16'h525F	;
				14'b01100011100010: Data_out <= 16'h5255	;
				14'b01100011100011: Data_out <= 16'h524C	;
				14'b01100011100100: Data_out <= 16'h5242	;
				14'b01100011100101: Data_out <= 16'h5238	;
				14'b01100011100110: Data_out <= 16'h522F	;
				14'b01100011100111: Data_out <= 16'h5225	;
				14'b01100011101000: Data_out <= 16'h521C	;
				14'b01100011101001: Data_out <= 16'h5212	;
				14'b01100011101010: Data_out <= 16'h5208	;
				14'b01100011101011: Data_out <= 16'h51FF	;
				14'b01100011101100: Data_out <= 16'h51F5	;
				14'b01100011101101: Data_out <= 16'h51EB	;
				14'b01100011101110: Data_out <= 16'h51E2	;
				14'b01100011101111: Data_out <= 16'h51D8	;
				14'b01100011110000: Data_out <= 16'h51CE	;
				14'b01100011110001: Data_out <= 16'h51C5	;
				14'b01100011110010: Data_out <= 16'h51BB	;
				14'b01100011110011: Data_out <= 16'h51B1	;
				14'b01100011110100: Data_out <= 16'h51A8	;
				14'b01100011110101: Data_out <= 16'h519E	;
				14'b01100011110110: Data_out <= 16'h5194	;
				14'b01100011110111: Data_out <= 16'h518B	;
				14'b01100011111000: Data_out <= 16'h5181	;
				14'b01100011111001: Data_out <= 16'h5177	;
				14'b01100011111010: Data_out <= 16'h516D	;
				14'b01100011111011: Data_out <= 16'h5164	;
				14'b01100011111100: Data_out <= 16'h515A	;
				14'b01100011111101: Data_out <= 16'h5150	;
				14'b01100011111110: Data_out <= 16'h5147	;
				14'b01100011111111: Data_out <= 16'h513D	;
				14'b01100100000000: Data_out <= 16'h5133	;
				14'b01100100000001: Data_out <= 16'h512A	;
				14'b01100100000010: Data_out <= 16'h5120	;
				14'b01100100000011: Data_out <= 16'h5116	;
				14'b01100100000100: Data_out <= 16'h510C	;
				14'b01100100000101: Data_out <= 16'h5103	;
				14'b01100100000110: Data_out <= 16'h50F9	;
				14'b01100100000111: Data_out <= 16'h50EF	;
				14'b01100100001000: Data_out <= 16'h50E5	;
				14'b01100100001001: Data_out <= 16'h50DC	;
				14'b01100100001010: Data_out <= 16'h50D2	;
				14'b01100100001011: Data_out <= 16'h50C8	;
				14'b01100100001100: Data_out <= 16'h50BE	;
				14'b01100100001101: Data_out <= 16'h50B5	;
				14'b01100100001110: Data_out <= 16'h50AB	;
				14'b01100100001111: Data_out <= 16'h50A1	;
				14'b01100100010000: Data_out <= 16'h5097	;
				14'b01100100010001: Data_out <= 16'h508E	;
				14'b01100100010010: Data_out <= 16'h5084	;
				14'b01100100010011: Data_out <= 16'h507A	;
				14'b01100100010100: Data_out <= 16'h5070	;
				14'b01100100010101: Data_out <= 16'h5067	;
				14'b01100100010110: Data_out <= 16'h505D	;
				14'b01100100010111: Data_out <= 16'h5053	;
				14'b01100100011000: Data_out <= 16'h5049	;
				14'b01100100011001: Data_out <= 16'h503F	;
				14'b01100100011010: Data_out <= 16'h5036	;
				14'b01100100011011: Data_out <= 16'h502C	;
				14'b01100100011100: Data_out <= 16'h5022	;
				14'b01100100011101: Data_out <= 16'h5018	;
				14'b01100100011110: Data_out <= 16'h500E	;
				14'b01100100011111: Data_out <= 16'h5005	;
				14'b01100100100000: Data_out <= 16'h4FFB	;
				14'b01100100100001: Data_out <= 16'h4FF1	;
				14'b01100100100010: Data_out <= 16'h4FE7	;
				14'b01100100100011: Data_out <= 16'h4FDD	;
				14'b01100100100100: Data_out <= 16'h4FD4	;
				14'b01100100100101: Data_out <= 16'h4FCA	;
				14'b01100100100110: Data_out <= 16'h4FC0	;
				14'b01100100100111: Data_out <= 16'h4FB6	;
				14'b01100100101000: Data_out <= 16'h4FAC	;
				14'b01100100101001: Data_out <= 16'h4FA2	;
				14'b01100100101010: Data_out <= 16'h4F99	;
				14'b01100100101011: Data_out <= 16'h4F8F	;
				14'b01100100101100: Data_out <= 16'h4F85	;
				14'b01100100101101: Data_out <= 16'h4F7B	;
				14'b01100100101110: Data_out <= 16'h4F71	;
				14'b01100100101111: Data_out <= 16'h4F67	;
				14'b01100100110000: Data_out <= 16'h4F5E	;
				14'b01100100110001: Data_out <= 16'h4F54	;
				14'b01100100110010: Data_out <= 16'h4F4A	;
				14'b01100100110011: Data_out <= 16'h4F40	;
				14'b01100100110100: Data_out <= 16'h4F36	;
				14'b01100100110101: Data_out <= 16'h4F2C	;
				14'b01100100110110: Data_out <= 16'h4F22	;
				14'b01100100110111: Data_out <= 16'h4F18	;
				14'b01100100111000: Data_out <= 16'h4F0F	;
				14'b01100100111001: Data_out <= 16'h4F05	;
				14'b01100100111010: Data_out <= 16'h4EFB	;
				14'b01100100111011: Data_out <= 16'h4EF1	;
				14'b01100100111100: Data_out <= 16'h4EE7	;
				14'b01100100111101: Data_out <= 16'h4EDD	;
				14'b01100100111110: Data_out <= 16'h4ED3	;
				14'b01100100111111: Data_out <= 16'h4EC9	;
				14'b01100101000000: Data_out <= 16'h4EBF	;
				14'b01100101000001: Data_out <= 16'h4EB5	;
				14'b01100101000010: Data_out <= 16'h4EAC	;
				14'b01100101000011: Data_out <= 16'h4EA2	;
				14'b01100101000100: Data_out <= 16'h4E98	;
				14'b01100101000101: Data_out <= 16'h4E8E	;
				14'b01100101000110: Data_out <= 16'h4E84	;
				14'b01100101000111: Data_out <= 16'h4E7A	;
				14'b01100101001000: Data_out <= 16'h4E70	;
				14'b01100101001001: Data_out <= 16'h4E66	;
				14'b01100101001010: Data_out <= 16'h4E5C	;
				14'b01100101001011: Data_out <= 16'h4E52	;
				14'b01100101001100: Data_out <= 16'h4E48	;
				14'b01100101001101: Data_out <= 16'h4E3E	;
				14'b01100101001110: Data_out <= 16'h4E34	;
				14'b01100101001111: Data_out <= 16'h4E2A	;
				14'b01100101010000: Data_out <= 16'h4E21	;
				14'b01100101010001: Data_out <= 16'h4E17	;
				14'b01100101010010: Data_out <= 16'h4E0D	;
				14'b01100101010011: Data_out <= 16'h4E03	;
				14'b01100101010100: Data_out <= 16'h4DF9	;
				14'b01100101010101: Data_out <= 16'h4DEF	;
				14'b01100101010110: Data_out <= 16'h4DE5	;
				14'b01100101010111: Data_out <= 16'h4DDB	;
				14'b01100101011000: Data_out <= 16'h4DD1	;
				14'b01100101011001: Data_out <= 16'h4DC7	;
				14'b01100101011010: Data_out <= 16'h4DBD	;
				14'b01100101011011: Data_out <= 16'h4DB3	;
				14'b01100101011100: Data_out <= 16'h4DA9	;
				14'b01100101011101: Data_out <= 16'h4D9F	;
				14'b01100101011110: Data_out <= 16'h4D95	;
				14'b01100101011111: Data_out <= 16'h4D8B	;
				14'b01100101100000: Data_out <= 16'h4D81	;
				14'b01100101100001: Data_out <= 16'h4D77	;
				14'b01100101100010: Data_out <= 16'h4D6D	;
				14'b01100101100011: Data_out <= 16'h4D63	;
				14'b01100101100100: Data_out <= 16'h4D59	;
				14'b01100101100101: Data_out <= 16'h4D4F	;
				14'b01100101100110: Data_out <= 16'h4D45	;
				14'b01100101100111: Data_out <= 16'h4D3B	;
				14'b01100101101000: Data_out <= 16'h4D31	;
				14'b01100101101001: Data_out <= 16'h4D27	;
				14'b01100101101010: Data_out <= 16'h4D1D	;
				14'b01100101101011: Data_out <= 16'h4D13	;
				14'b01100101101100: Data_out <= 16'h4D09	;
				14'b01100101101101: Data_out <= 16'h4CFF	;
				14'b01100101101110: Data_out <= 16'h4CF5	;
				14'b01100101101111: Data_out <= 16'h4CEB	;
				14'b01100101110000: Data_out <= 16'h4CE1	;
				14'b01100101110001: Data_out <= 16'h4CD6	;
				14'b01100101110010: Data_out <= 16'h4CCC	;
				14'b01100101110011: Data_out <= 16'h4CC2	;
				14'b01100101110100: Data_out <= 16'h4CB8	;
				14'b01100101110101: Data_out <= 16'h4CAE	;
				14'b01100101110110: Data_out <= 16'h4CA4	;
				14'b01100101110111: Data_out <= 16'h4C9A	;
				14'b01100101111000: Data_out <= 16'h4C90	;
				14'b01100101111001: Data_out <= 16'h4C86	;
				14'b01100101111010: Data_out <= 16'h4C7C	;
				14'b01100101111011: Data_out <= 16'h4C72	;
				14'b01100101111100: Data_out <= 16'h4C68	;
				14'b01100101111101: Data_out <= 16'h4C5E	;
				14'b01100101111110: Data_out <= 16'h4C54	;
				14'b01100101111111: Data_out <= 16'h4C49	;
				14'b01100110000000: Data_out <= 16'h4C3F	;
				14'b01100110000001: Data_out <= 16'h4C35	;
				14'b01100110000010: Data_out <= 16'h4C2B	;
				14'b01100110000011: Data_out <= 16'h4C21	;
				14'b01100110000100: Data_out <= 16'h4C17	;
				14'b01100110000101: Data_out <= 16'h4C0D	;
				14'b01100110000110: Data_out <= 16'h4C03	;
				14'b01100110000111: Data_out <= 16'h4BF9	;
				14'b01100110001000: Data_out <= 16'h4BEF	;
				14'b01100110001001: Data_out <= 16'h4BE4	;
				14'b01100110001010: Data_out <= 16'h4BDA	;
				14'b01100110001011: Data_out <= 16'h4BD0	;
				14'b01100110001100: Data_out <= 16'h4BC6	;
				14'b01100110001101: Data_out <= 16'h4BBC	;
				14'b01100110001110: Data_out <= 16'h4BB2	;
				14'b01100110001111: Data_out <= 16'h4BA8	;
				14'b01100110010000: Data_out <= 16'h4B9E	;
				14'b01100110010001: Data_out <= 16'h4B93	;
				14'b01100110010010: Data_out <= 16'h4B89	;
				14'b01100110010011: Data_out <= 16'h4B7F	;
				14'b01100110010100: Data_out <= 16'h4B75	;
				14'b01100110010101: Data_out <= 16'h4B6B	;
				14'b01100110010110: Data_out <= 16'h4B61	;
				14'b01100110010111: Data_out <= 16'h4B56	;
				14'b01100110011000: Data_out <= 16'h4B4C	;
				14'b01100110011001: Data_out <= 16'h4B42	;
				14'b01100110011010: Data_out <= 16'h4B38	;
				14'b01100110011011: Data_out <= 16'h4B2E	;
				14'b01100110011100: Data_out <= 16'h4B24	;
				14'b01100110011101: Data_out <= 16'h4B19	;
				14'b01100110011110: Data_out <= 16'h4B0F	;
				14'b01100110011111: Data_out <= 16'h4B05	;
				14'b01100110100000: Data_out <= 16'h4AFB	;
				14'b01100110100001: Data_out <= 16'h4AF1	;
				14'b01100110100010: Data_out <= 16'h4AE7	;
				14'b01100110100011: Data_out <= 16'h4ADC	;
				14'b01100110100100: Data_out <= 16'h4AD2	;
				14'b01100110100101: Data_out <= 16'h4AC8	;
				14'b01100110100110: Data_out <= 16'h4ABE	;
				14'b01100110100111: Data_out <= 16'h4AB4	;
				14'b01100110101000: Data_out <= 16'h4AA9	;
				14'b01100110101001: Data_out <= 16'h4A9F	;
				14'b01100110101010: Data_out <= 16'h4A95	;
				14'b01100110101011: Data_out <= 16'h4A8B	;
				14'b01100110101100: Data_out <= 16'h4A81	;
				14'b01100110101101: Data_out <= 16'h4A76	;
				14'b01100110101110: Data_out <= 16'h4A6C	;
				14'b01100110101111: Data_out <= 16'h4A62	;
				14'b01100110110000: Data_out <= 16'h4A58	;
				14'b01100110110001: Data_out <= 16'h4A4D	;
				14'b01100110110010: Data_out <= 16'h4A43	;
				14'b01100110110011: Data_out <= 16'h4A39	;
				14'b01100110110100: Data_out <= 16'h4A2F	;
				14'b01100110110101: Data_out <= 16'h4A24	;
				14'b01100110110110: Data_out <= 16'h4A1A	;
				14'b01100110110111: Data_out <= 16'h4A10	;
				14'b01100110111000: Data_out <= 16'h4A06	;
				14'b01100110111001: Data_out <= 16'h49FB	;
				14'b01100110111010: Data_out <= 16'h49F1	;
				14'b01100110111011: Data_out <= 16'h49E7	;
				14'b01100110111100: Data_out <= 16'h49DD	;
				14'b01100110111101: Data_out <= 16'h49D2	;
				14'b01100110111110: Data_out <= 16'h49C8	;
				14'b01100110111111: Data_out <= 16'h49BE	;
				14'b01100111000000: Data_out <= 16'h49B4	;
				14'b01100111000001: Data_out <= 16'h49A9	;
				14'b01100111000010: Data_out <= 16'h499F	;
				14'b01100111000011: Data_out <= 16'h4995	;
				14'b01100111000100: Data_out <= 16'h498A	;
				14'b01100111000101: Data_out <= 16'h4980	;
				14'b01100111000110: Data_out <= 16'h4976	;
				14'b01100111000111: Data_out <= 16'h496C	;
				14'b01100111001000: Data_out <= 16'h4961	;
				14'b01100111001001: Data_out <= 16'h4957	;
				14'b01100111001010: Data_out <= 16'h494D	;
				14'b01100111001011: Data_out <= 16'h4942	;
				14'b01100111001100: Data_out <= 16'h4938	;
				14'b01100111001101: Data_out <= 16'h492E	;
				14'b01100111001110: Data_out <= 16'h4924	;
				14'b01100111001111: Data_out <= 16'h4919	;
				14'b01100111010000: Data_out <= 16'h490F	;
				14'b01100111010001: Data_out <= 16'h4905	;
				14'b01100111010010: Data_out <= 16'h48FA	;
				14'b01100111010011: Data_out <= 16'h48F0	;
				14'b01100111010100: Data_out <= 16'h48E6	;
				14'b01100111010101: Data_out <= 16'h48DB	;
				14'b01100111010110: Data_out <= 16'h48D1	;
				14'b01100111010111: Data_out <= 16'h48C7	;
				14'b01100111011000: Data_out <= 16'h48BC	;
				14'b01100111011001: Data_out <= 16'h48B2	;
				14'b01100111011010: Data_out <= 16'h48A8	;
				14'b01100111011011: Data_out <= 16'h489D	;
				14'b01100111011100: Data_out <= 16'h4893	;
				14'b01100111011101: Data_out <= 16'h4889	;
				14'b01100111011110: Data_out <= 16'h487E	;
				14'b01100111011111: Data_out <= 16'h4874	;
				14'b01100111100000: Data_out <= 16'h4869	;
				14'b01100111100001: Data_out <= 16'h485F	;
				14'b01100111100010: Data_out <= 16'h4855	;
				14'b01100111100011: Data_out <= 16'h484A	;
				14'b01100111100100: Data_out <= 16'h4840	;
				14'b01100111100101: Data_out <= 16'h4836	;
				14'b01100111100110: Data_out <= 16'h482B	;
				14'b01100111100111: Data_out <= 16'h4821	;
				14'b01100111101000: Data_out <= 16'h4816	;
				14'b01100111101001: Data_out <= 16'h480C	;
				14'b01100111101010: Data_out <= 16'h4802	;
				14'b01100111101011: Data_out <= 16'h47F7	;
				14'b01100111101100: Data_out <= 16'h47ED	;
				14'b01100111101101: Data_out <= 16'h47E3	;
				14'b01100111101110: Data_out <= 16'h47D8	;
				14'b01100111101111: Data_out <= 16'h47CE	;
				14'b01100111110000: Data_out <= 16'h47C3	;
				14'b01100111110001: Data_out <= 16'h47B9	;
				14'b01100111110010: Data_out <= 16'h47AE	;
				14'b01100111110011: Data_out <= 16'h47A4	;
				14'b01100111110100: Data_out <= 16'h479A	;
				14'b01100111110101: Data_out <= 16'h478F	;
				14'b01100111110110: Data_out <= 16'h4785	;
				14'b01100111110111: Data_out <= 16'h477A	;
				14'b01100111111000: Data_out <= 16'h4770	;
				14'b01100111111001: Data_out <= 16'h4766	;
				14'b01100111111010: Data_out <= 16'h475B	;
				14'b01100111111011: Data_out <= 16'h4751	;
				14'b01100111111100: Data_out <= 16'h4746	;
				14'b01100111111101: Data_out <= 16'h473C	;
				14'b01100111111110: Data_out <= 16'h4731	;
				14'b01100111111111: Data_out <= 16'h4727	;
				14'b01101000000000: Data_out <= 16'h471C	;
				14'b01101000000001: Data_out <= 16'h4712	;
				14'b01101000000010: Data_out <= 16'h4708	;
				14'b01101000000011: Data_out <= 16'h46FD	;
				14'b01101000000100: Data_out <= 16'h46F3	;
				14'b01101000000101: Data_out <= 16'h46E8	;
				14'b01101000000110: Data_out <= 16'h46DE	;
				14'b01101000000111: Data_out <= 16'h46D3	;
				14'b01101000001000: Data_out <= 16'h46C9	;
				14'b01101000001001: Data_out <= 16'h46BE	;
				14'b01101000001010: Data_out <= 16'h46B4	;
				14'b01101000001011: Data_out <= 16'h46A9	;
				14'b01101000001100: Data_out <= 16'h469F	;
				14'b01101000001101: Data_out <= 16'h4694	;
				14'b01101000001110: Data_out <= 16'h468A	;
				14'b01101000001111: Data_out <= 16'h467F	;
				14'b01101000010000: Data_out <= 16'h4675	;
				14'b01101000010001: Data_out <= 16'h466A	;
				14'b01101000010010: Data_out <= 16'h4660	;
				14'b01101000010011: Data_out <= 16'h4655	;
				14'b01101000010100: Data_out <= 16'h464B	;
				14'b01101000010101: Data_out <= 16'h4640	;
				14'b01101000010110: Data_out <= 16'h4636	;
				14'b01101000010111: Data_out <= 16'h462B	;
				14'b01101000011000: Data_out <= 16'h4621	;
				14'b01101000011001: Data_out <= 16'h4616	;
				14'b01101000011010: Data_out <= 16'h460C	;
				14'b01101000011011: Data_out <= 16'h4601	;
				14'b01101000011100: Data_out <= 16'h45F7	;
				14'b01101000011101: Data_out <= 16'h45EC	;
				14'b01101000011110: Data_out <= 16'h45E2	;
				14'b01101000011111: Data_out <= 16'h45D7	;
				14'b01101000100000: Data_out <= 16'h45CD	;
				14'b01101000100001: Data_out <= 16'h45C2	;
				14'b01101000100010: Data_out <= 16'h45B8	;
				14'b01101000100011: Data_out <= 16'h45AD	;
				14'b01101000100100: Data_out <= 16'h45A3	;
				14'b01101000100101: Data_out <= 16'h4598	;
				14'b01101000100110: Data_out <= 16'h458E	;
				14'b01101000100111: Data_out <= 16'h4583	;
				14'b01101000101000: Data_out <= 16'h4578	;
				14'b01101000101001: Data_out <= 16'h456E	;
				14'b01101000101010: Data_out <= 16'h4563	;
				14'b01101000101011: Data_out <= 16'h4559	;
				14'b01101000101100: Data_out <= 16'h454E	;
				14'b01101000101101: Data_out <= 16'h4544	;
				14'b01101000101110: Data_out <= 16'h4539	;
				14'b01101000101111: Data_out <= 16'h452E	;
				14'b01101000110000: Data_out <= 16'h4524	;
				14'b01101000110001: Data_out <= 16'h4519	;
				14'b01101000110010: Data_out <= 16'h450F	;
				14'b01101000110011: Data_out <= 16'h4504	;
				14'b01101000110100: Data_out <= 16'h44FA	;
				14'b01101000110101: Data_out <= 16'h44EF	;
				14'b01101000110110: Data_out <= 16'h44E4	;
				14'b01101000110111: Data_out <= 16'h44DA	;
				14'b01101000111000: Data_out <= 16'h44CF	;
				14'b01101000111001: Data_out <= 16'h44C5	;
				14'b01101000111010: Data_out <= 16'h44BA	;
				14'b01101000111011: Data_out <= 16'h44AF	;
				14'b01101000111100: Data_out <= 16'h44A5	;
				14'b01101000111101: Data_out <= 16'h449A	;
				14'b01101000111110: Data_out <= 16'h4490	;
				14'b01101000111111: Data_out <= 16'h4485	;
				14'b01101001000000: Data_out <= 16'h447A	;
				14'b01101001000001: Data_out <= 16'h4470	;
				14'b01101001000010: Data_out <= 16'h4465	;
				14'b01101001000011: Data_out <= 16'h445B	;
				14'b01101001000100: Data_out <= 16'h4450	;
				14'b01101001000101: Data_out <= 16'h4445	;
				14'b01101001000110: Data_out <= 16'h443B	;
				14'b01101001000111: Data_out <= 16'h4430	;
				14'b01101001001000: Data_out <= 16'h4425	;
				14'b01101001001001: Data_out <= 16'h441B	;
				14'b01101001001010: Data_out <= 16'h4410	;
				14'b01101001001011: Data_out <= 16'h4405	;
				14'b01101001001100: Data_out <= 16'h43FB	;
				14'b01101001001101: Data_out <= 16'h43F0	;
				14'b01101001001110: Data_out <= 16'h43E5	;
				14'b01101001001111: Data_out <= 16'h43DB	;
				14'b01101001010000: Data_out <= 16'h43D0	;
				14'b01101001010001: Data_out <= 16'h43C6	;
				14'b01101001010010: Data_out <= 16'h43BB	;
				14'b01101001010011: Data_out <= 16'h43B0	;
				14'b01101001010100: Data_out <= 16'h43A6	;
				14'b01101001010101: Data_out <= 16'h439B	;
				14'b01101001010110: Data_out <= 16'h4390	;
				14'b01101001010111: Data_out <= 16'h4386	;
				14'b01101001011000: Data_out <= 16'h437B	;
				14'b01101001011001: Data_out <= 16'h4370	;
				14'b01101001011010: Data_out <= 16'h4365	;
				14'b01101001011011: Data_out <= 16'h435B	;
				14'b01101001011100: Data_out <= 16'h4350	;
				14'b01101001011101: Data_out <= 16'h4345	;
				14'b01101001011110: Data_out <= 16'h433B	;
				14'b01101001011111: Data_out <= 16'h4330	;
				14'b01101001100000: Data_out <= 16'h4325	;
				14'b01101001100001: Data_out <= 16'h431B	;
				14'b01101001100010: Data_out <= 16'h4310	;
				14'b01101001100011: Data_out <= 16'h4305	;
				14'b01101001100100: Data_out <= 16'h42FB	;
				14'b01101001100101: Data_out <= 16'h42F0	;
				14'b01101001100110: Data_out <= 16'h42E5	;
				14'b01101001100111: Data_out <= 16'h42DA	;
				14'b01101001101000: Data_out <= 16'h42D0	;
				14'b01101001101001: Data_out <= 16'h42C5	;
				14'b01101001101010: Data_out <= 16'h42BA	;
				14'b01101001101011: Data_out <= 16'h42AF	;
				14'b01101001101100: Data_out <= 16'h42A5	;
				14'b01101001101101: Data_out <= 16'h429A	;
				14'b01101001101110: Data_out <= 16'h428F	;
				14'b01101001101111: Data_out <= 16'h4285	;
				14'b01101001110000: Data_out <= 16'h427A	;
				14'b01101001110001: Data_out <= 16'h426F	;
				14'b01101001110010: Data_out <= 16'h4264	;
				14'b01101001110011: Data_out <= 16'h425A	;
				14'b01101001110100: Data_out <= 16'h424F	;
				14'b01101001110101: Data_out <= 16'h4244	;
				14'b01101001110110: Data_out <= 16'h4239	;
				14'b01101001110111: Data_out <= 16'h422F	;
				14'b01101001111000: Data_out <= 16'h4224	;
				14'b01101001111001: Data_out <= 16'h4219	;
				14'b01101001111010: Data_out <= 16'h420E	;
				14'b01101001111011: Data_out <= 16'h4204	;
				14'b01101001111100: Data_out <= 16'h41F9	;
				14'b01101001111101: Data_out <= 16'h41EE	;
				14'b01101001111110: Data_out <= 16'h41E3	;
				14'b01101001111111: Data_out <= 16'h41D8	;
				14'b01101010000000: Data_out <= 16'h41CE	;
				14'b01101010000001: Data_out <= 16'h41C3	;
				14'b01101010000010: Data_out <= 16'h41B8	;
				14'b01101010000011: Data_out <= 16'h41AD	;
				14'b01101010000100: Data_out <= 16'h41A3	;
				14'b01101010000101: Data_out <= 16'h4198	;
				14'b01101010000110: Data_out <= 16'h418D	;
				14'b01101010000111: Data_out <= 16'h4182	;
				14'b01101010001000: Data_out <= 16'h4177	;
				14'b01101010001001: Data_out <= 16'h416D	;
				14'b01101010001010: Data_out <= 16'h4162	;
				14'b01101010001011: Data_out <= 16'h4157	;
				14'b01101010001100: Data_out <= 16'h414C	;
				14'b01101010001101: Data_out <= 16'h4141	;
				14'b01101010001110: Data_out <= 16'h4137	;
				14'b01101010001111: Data_out <= 16'h412C	;
				14'b01101010010000: Data_out <= 16'h4121	;
				14'b01101010010001: Data_out <= 16'h4116	;
				14'b01101010010010: Data_out <= 16'h410B	;
				14'b01101010010011: Data_out <= 16'h4100	;
				14'b01101010010100: Data_out <= 16'h40F6	;
				14'b01101010010101: Data_out <= 16'h40EB	;
				14'b01101010010110: Data_out <= 16'h40E0	;
				14'b01101010010111: Data_out <= 16'h40D5	;
				14'b01101010011000: Data_out <= 16'h40CA	;
				14'b01101010011001: Data_out <= 16'h40BF	;
				14'b01101010011010: Data_out <= 16'h40B5	;
				14'b01101010011011: Data_out <= 16'h40AA	;
				14'b01101010011100: Data_out <= 16'h409F	;
				14'b01101010011101: Data_out <= 16'h4094	;
				14'b01101010011110: Data_out <= 16'h4089	;
				14'b01101010011111: Data_out <= 16'h407E	;
				14'b01101010100000: Data_out <= 16'h4074	;
				14'b01101010100001: Data_out <= 16'h4069	;
				14'b01101010100010: Data_out <= 16'h405E	;
				14'b01101010100011: Data_out <= 16'h4053	;
				14'b01101010100100: Data_out <= 16'h4048	;
				14'b01101010100101: Data_out <= 16'h403D	;
				14'b01101010100110: Data_out <= 16'h4032	;
				14'b01101010100111: Data_out <= 16'h4027	;
				14'b01101010101000: Data_out <= 16'h401D	;
				14'b01101010101001: Data_out <= 16'h4012	;
				14'b01101010101010: Data_out <= 16'h4007	;
				14'b01101010101011: Data_out <= 16'h3FFC	;
				14'b01101010101100: Data_out <= 16'h3FF1	;
				14'b01101010101101: Data_out <= 16'h3FE6	;
				14'b01101010101110: Data_out <= 16'h3FDB	;
				14'b01101010101111: Data_out <= 16'h3FD0	;
				14'b01101010110000: Data_out <= 16'h3FC6	;
				14'b01101010110001: Data_out <= 16'h3FBB	;
				14'b01101010110010: Data_out <= 16'h3FB0	;
				14'b01101010110011: Data_out <= 16'h3FA5	;
				14'b01101010110100: Data_out <= 16'h3F9A	;
				14'b01101010110101: Data_out <= 16'h3F8F	;
				14'b01101010110110: Data_out <= 16'h3F84	;
				14'b01101010110111: Data_out <= 16'h3F79	;
				14'b01101010111000: Data_out <= 16'h3F6E	;
				14'b01101010111001: Data_out <= 16'h3F63	;
				14'b01101010111010: Data_out <= 16'h3F58	;
				14'b01101010111011: Data_out <= 16'h3F4E	;
				14'b01101010111100: Data_out <= 16'h3F43	;
				14'b01101010111101: Data_out <= 16'h3F38	;
				14'b01101010111110: Data_out <= 16'h3F2D	;
				14'b01101010111111: Data_out <= 16'h3F22	;
				14'b01101011000000: Data_out <= 16'h3F17	;
				14'b01101011000001: Data_out <= 16'h3F0C	;
				14'b01101011000010: Data_out <= 16'h3F01	;
				14'b01101011000011: Data_out <= 16'h3EF6	;
				14'b01101011000100: Data_out <= 16'h3EEB	;
				14'b01101011000101: Data_out <= 16'h3EE0	;
				14'b01101011000110: Data_out <= 16'h3ED5	;
				14'b01101011000111: Data_out <= 16'h3ECA	;
				14'b01101011001000: Data_out <= 16'h3EBF	;
				14'b01101011001001: Data_out <= 16'h3EB4	;
				14'b01101011001010: Data_out <= 16'h3EA9	;
				14'b01101011001011: Data_out <= 16'h3E9E	;
				14'b01101011001100: Data_out <= 16'h3E94	;
				14'b01101011001101: Data_out <= 16'h3E89	;
				14'b01101011001110: Data_out <= 16'h3E7E	;
				14'b01101011001111: Data_out <= 16'h3E73	;
				14'b01101011010000: Data_out <= 16'h3E68	;
				14'b01101011010001: Data_out <= 16'h3E5D	;
				14'b01101011010010: Data_out <= 16'h3E52	;
				14'b01101011010011: Data_out <= 16'h3E47	;
				14'b01101011010100: Data_out <= 16'h3E3C	;
				14'b01101011010101: Data_out <= 16'h3E31	;
				14'b01101011010110: Data_out <= 16'h3E26	;
				14'b01101011010111: Data_out <= 16'h3E1B	;
				14'b01101011011000: Data_out <= 16'h3E10	;
				14'b01101011011001: Data_out <= 16'h3E05	;
				14'b01101011011010: Data_out <= 16'h3DFA	;
				14'b01101011011011: Data_out <= 16'h3DEF	;
				14'b01101011011100: Data_out <= 16'h3DE4	;
				14'b01101011011101: Data_out <= 16'h3DD9	;
				14'b01101011011110: Data_out <= 16'h3DCE	;
				14'b01101011011111: Data_out <= 16'h3DC3	;
				14'b01101011100000: Data_out <= 16'h3DB8	;
				14'b01101011100001: Data_out <= 16'h3DAD	;
				14'b01101011100010: Data_out <= 16'h3DA2	;
				14'b01101011100011: Data_out <= 16'h3D97	;
				14'b01101011100100: Data_out <= 16'h3D8C	;
				14'b01101011100101: Data_out <= 16'h3D81	;
				14'b01101011100110: Data_out <= 16'h3D76	;
				14'b01101011100111: Data_out <= 16'h3D6B	;
				14'b01101011101000: Data_out <= 16'h3D60	;
				14'b01101011101001: Data_out <= 16'h3D55	;
				14'b01101011101010: Data_out <= 16'h3D4A	;
				14'b01101011101011: Data_out <= 16'h3D3F	;
				14'b01101011101100: Data_out <= 16'h3D34	;
				14'b01101011101101: Data_out <= 16'h3D29	;
				14'b01101011101110: Data_out <= 16'h3D1D	;
				14'b01101011101111: Data_out <= 16'h3D12	;
				14'b01101011110000: Data_out <= 16'h3D07	;
				14'b01101011110001: Data_out <= 16'h3CFC	;
				14'b01101011110010: Data_out <= 16'h3CF1	;
				14'b01101011110011: Data_out <= 16'h3CE6	;
				14'b01101011110100: Data_out <= 16'h3CDB	;
				14'b01101011110101: Data_out <= 16'h3CD0	;
				14'b01101011110110: Data_out <= 16'h3CC5	;
				14'b01101011110111: Data_out <= 16'h3CBA	;
				14'b01101011111000: Data_out <= 16'h3CAF	;
				14'b01101011111001: Data_out <= 16'h3CA4	;
				14'b01101011111010: Data_out <= 16'h3C99	;
				14'b01101011111011: Data_out <= 16'h3C8E	;
				14'b01101011111100: Data_out <= 16'h3C83	;
				14'b01101011111101: Data_out <= 16'h3C78	;
				14'b01101011111110: Data_out <= 16'h3C6D	;
				14'b01101011111111: Data_out <= 16'h3C61	;
				14'b01101100000000: Data_out <= 16'h3C56	;
				14'b01101100000001: Data_out <= 16'h3C4B	;
				14'b01101100000010: Data_out <= 16'h3C40	;
				14'b01101100000011: Data_out <= 16'h3C35	;
				14'b01101100000100: Data_out <= 16'h3C2A	;
				14'b01101100000101: Data_out <= 16'h3C1F	;
				14'b01101100000110: Data_out <= 16'h3C14	;
				14'b01101100000111: Data_out <= 16'h3C09	;
				14'b01101100001000: Data_out <= 16'h3BFE	;
				14'b01101100001001: Data_out <= 16'h3BF3	;
				14'b01101100001010: Data_out <= 16'h3BE7	;
				14'b01101100001011: Data_out <= 16'h3BDC	;
				14'b01101100001100: Data_out <= 16'h3BD1	;
				14'b01101100001101: Data_out <= 16'h3BC6	;
				14'b01101100001110: Data_out <= 16'h3BBB	;
				14'b01101100001111: Data_out <= 16'h3BB0	;
				14'b01101100010000: Data_out <= 16'h3BA5	;
				14'b01101100010001: Data_out <= 16'h3B9A	;
				14'b01101100010010: Data_out <= 16'h3B8F	;
				14'b01101100010011: Data_out <= 16'h3B83	;
				14'b01101100010100: Data_out <= 16'h3B78	;
				14'b01101100010101: Data_out <= 16'h3B6D	;
				14'b01101100010110: Data_out <= 16'h3B62	;
				14'b01101100010111: Data_out <= 16'h3B57	;
				14'b01101100011000: Data_out <= 16'h3B4C	;
				14'b01101100011001: Data_out <= 16'h3B41	;
				14'b01101100011010: Data_out <= 16'h3B35	;
				14'b01101100011011: Data_out <= 16'h3B2A	;
				14'b01101100011100: Data_out <= 16'h3B1F	;
				14'b01101100011101: Data_out <= 16'h3B14	;
				14'b01101100011110: Data_out <= 16'h3B09	;
				14'b01101100011111: Data_out <= 16'h3AFE	;
				14'b01101100100000: Data_out <= 16'h3AF3	;
				14'b01101100100001: Data_out <= 16'h3AE7	;
				14'b01101100100010: Data_out <= 16'h3ADC	;
				14'b01101100100011: Data_out <= 16'h3AD1	;
				14'b01101100100100: Data_out <= 16'h3AC6	;
				14'b01101100100101: Data_out <= 16'h3ABB	;
				14'b01101100100110: Data_out <= 16'h3AB0	;
				14'b01101100100111: Data_out <= 16'h3AA4	;
				14'b01101100101000: Data_out <= 16'h3A99	;
				14'b01101100101001: Data_out <= 16'h3A8E	;
				14'b01101100101010: Data_out <= 16'h3A83	;
				14'b01101100101011: Data_out <= 16'h3A78	;
				14'b01101100101100: Data_out <= 16'h3A6D	;
				14'b01101100101101: Data_out <= 16'h3A61	;
				14'b01101100101110: Data_out <= 16'h3A56	;
				14'b01101100101111: Data_out <= 16'h3A4B	;
				14'b01101100110000: Data_out <= 16'h3A40	;
				14'b01101100110001: Data_out <= 16'h3A35	;
				14'b01101100110010: Data_out <= 16'h3A29	;
				14'b01101100110011: Data_out <= 16'h3A1E	;
				14'b01101100110100: Data_out <= 16'h3A13	;
				14'b01101100110101: Data_out <= 16'h3A08	;
				14'b01101100110110: Data_out <= 16'h39FD	;
				14'b01101100110111: Data_out <= 16'h39F1	;
				14'b01101100111000: Data_out <= 16'h39E6	;
				14'b01101100111001: Data_out <= 16'h39DB	;
				14'b01101100111010: Data_out <= 16'h39D0	;
				14'b01101100111011: Data_out <= 16'h39C5	;
				14'b01101100111100: Data_out <= 16'h39B9	;
				14'b01101100111101: Data_out <= 16'h39AE	;
				14'b01101100111110: Data_out <= 16'h39A3	;
				14'b01101100111111: Data_out <= 16'h3998	;
				14'b01101101000000: Data_out <= 16'h398D	;
				14'b01101101000001: Data_out <= 16'h3981	;
				14'b01101101000010: Data_out <= 16'h3976	;
				14'b01101101000011: Data_out <= 16'h396B	;
				14'b01101101000100: Data_out <= 16'h3960	;
				14'b01101101000101: Data_out <= 16'h3954	;
				14'b01101101000110: Data_out <= 16'h3949	;
				14'b01101101000111: Data_out <= 16'h393E	;
				14'b01101101001000: Data_out <= 16'h3933	;
				14'b01101101001001: Data_out <= 16'h3927	;
				14'b01101101001010: Data_out <= 16'h391C	;
				14'b01101101001011: Data_out <= 16'h3911	;
				14'b01101101001100: Data_out <= 16'h3906	;
				14'b01101101001101: Data_out <= 16'h38FA	;
				14'b01101101001110: Data_out <= 16'h38EF	;
				14'b01101101001111: Data_out <= 16'h38E4	;
				14'b01101101010000: Data_out <= 16'h38D9	;
				14'b01101101010001: Data_out <= 16'h38CD	;
				14'b01101101010010: Data_out <= 16'h38C2	;
				14'b01101101010011: Data_out <= 16'h38B7	;
				14'b01101101010100: Data_out <= 16'h38AC	;
				14'b01101101010101: Data_out <= 16'h38A0	;
				14'b01101101010110: Data_out <= 16'h3895	;
				14'b01101101010111: Data_out <= 16'h388A	;
				14'b01101101011000: Data_out <= 16'h387F	;
				14'b01101101011001: Data_out <= 16'h3873	;
				14'b01101101011010: Data_out <= 16'h3868	;
				14'b01101101011011: Data_out <= 16'h385D	;
				14'b01101101011100: Data_out <= 16'h3851	;
				14'b01101101011101: Data_out <= 16'h3846	;
				14'b01101101011110: Data_out <= 16'h383B	;
				14'b01101101011111: Data_out <= 16'h3830	;
				14'b01101101100000: Data_out <= 16'h3824	;
				14'b01101101100001: Data_out <= 16'h3819	;
				14'b01101101100010: Data_out <= 16'h380E	;
				14'b01101101100011: Data_out <= 16'h3802	;
				14'b01101101100100: Data_out <= 16'h37F7	;
				14'b01101101100101: Data_out <= 16'h37EC	;
				14'b01101101100110: Data_out <= 16'h37E0	;
				14'b01101101100111: Data_out <= 16'h37D5	;
				14'b01101101101000: Data_out <= 16'h37CA	;
				14'b01101101101001: Data_out <= 16'h37BF	;
				14'b01101101101010: Data_out <= 16'h37B3	;
				14'b01101101101011: Data_out <= 16'h37A8	;
				14'b01101101101100: Data_out <= 16'h379D	;
				14'b01101101101101: Data_out <= 16'h3791	;
				14'b01101101101110: Data_out <= 16'h3786	;
				14'b01101101101111: Data_out <= 16'h377B	;
				14'b01101101110000: Data_out <= 16'h376F	;
				14'b01101101110001: Data_out <= 16'h3764	;
				14'b01101101110010: Data_out <= 16'h3759	;
				14'b01101101110011: Data_out <= 16'h374D	;
				14'b01101101110100: Data_out <= 16'h3742	;
				14'b01101101110101: Data_out <= 16'h3737	;
				14'b01101101110110: Data_out <= 16'h372B	;
				14'b01101101110111: Data_out <= 16'h3720	;
				14'b01101101111000: Data_out <= 16'h3715	;
				14'b01101101111001: Data_out <= 16'h3709	;
				14'b01101101111010: Data_out <= 16'h36FE	;
				14'b01101101111011: Data_out <= 16'h36F3	;
				14'b01101101111100: Data_out <= 16'h36E7	;
				14'b01101101111101: Data_out <= 16'h36DC	;
				14'b01101101111110: Data_out <= 16'h36D1	;
				14'b01101101111111: Data_out <= 16'h36C5	;
				14'b01101110000000: Data_out <= 16'h36BA	;
				14'b01101110000001: Data_out <= 16'h36AE	;
				14'b01101110000010: Data_out <= 16'h36A3	;
				14'b01101110000011: Data_out <= 16'h3698	;
				14'b01101110000100: Data_out <= 16'h368C	;
				14'b01101110000101: Data_out <= 16'h3681	;
				14'b01101110000110: Data_out <= 16'h3676	;
				14'b01101110000111: Data_out <= 16'h366A	;
				14'b01101110001000: Data_out <= 16'h365F	;
				14'b01101110001001: Data_out <= 16'h3653	;
				14'b01101110001010: Data_out <= 16'h3648	;
				14'b01101110001011: Data_out <= 16'h363D	;
				14'b01101110001100: Data_out <= 16'h3631	;
				14'b01101110001101: Data_out <= 16'h3626	;
				14'b01101110001110: Data_out <= 16'h361B	;
				14'b01101110001111: Data_out <= 16'h360F	;
				14'b01101110010000: Data_out <= 16'h3604	;
				14'b01101110010001: Data_out <= 16'h35F8	;
				14'b01101110010010: Data_out <= 16'h35ED	;
				14'b01101110010011: Data_out <= 16'h35E2	;
				14'b01101110010100: Data_out <= 16'h35D6	;
				14'b01101110010101: Data_out <= 16'h35CB	;
				14'b01101110010110: Data_out <= 16'h35BF	;
				14'b01101110010111: Data_out <= 16'h35B4	;
				14'b01101110011000: Data_out <= 16'h35A9	;
				14'b01101110011001: Data_out <= 16'h359D	;
				14'b01101110011010: Data_out <= 16'h3592	;
				14'b01101110011011: Data_out <= 16'h3586	;
				14'b01101110011100: Data_out <= 16'h357B	;
				14'b01101110011101: Data_out <= 16'h3570	;
				14'b01101110011110: Data_out <= 16'h3564	;
				14'b01101110011111: Data_out <= 16'h3559	;
				14'b01101110100000: Data_out <= 16'h354D	;
				14'b01101110100001: Data_out <= 16'h3542	;
				14'b01101110100010: Data_out <= 16'h3536	;
				14'b01101110100011: Data_out <= 16'h352B	;
				14'b01101110100100: Data_out <= 16'h3520	;
				14'b01101110100101: Data_out <= 16'h3514	;
				14'b01101110100110: Data_out <= 16'h3509	;
				14'b01101110100111: Data_out <= 16'h34FD	;
				14'b01101110101000: Data_out <= 16'h34F2	;
				14'b01101110101001: Data_out <= 16'h34E6	;
				14'b01101110101010: Data_out <= 16'h34DB	;
				14'b01101110101011: Data_out <= 16'h34CF	;
				14'b01101110101100: Data_out <= 16'h34C4	;
				14'b01101110101101: Data_out <= 16'h34B9	;
				14'b01101110101110: Data_out <= 16'h34AD	;
				14'b01101110101111: Data_out <= 16'h34A2	;
				14'b01101110110000: Data_out <= 16'h3496	;
				14'b01101110110001: Data_out <= 16'h348B	;
				14'b01101110110010: Data_out <= 16'h347F	;
				14'b01101110110011: Data_out <= 16'h3474	;
				14'b01101110110100: Data_out <= 16'h3468	;
				14'b01101110110101: Data_out <= 16'h345D	;
				14'b01101110110110: Data_out <= 16'h3451	;
				14'b01101110110111: Data_out <= 16'h3446	;
				14'b01101110111000: Data_out <= 16'h343A	;
				14'b01101110111001: Data_out <= 16'h342F	;
				14'b01101110111010: Data_out <= 16'h3424	;
				14'b01101110111011: Data_out <= 16'h3418	;
				14'b01101110111100: Data_out <= 16'h340D	;
				14'b01101110111101: Data_out <= 16'h3401	;
				14'b01101110111110: Data_out <= 16'h33F6	;
				14'b01101110111111: Data_out <= 16'h33EA	;
				14'b01101111000000: Data_out <= 16'h33DF	;
				14'b01101111000001: Data_out <= 16'h33D3	;
				14'b01101111000010: Data_out <= 16'h33C8	;
				14'b01101111000011: Data_out <= 16'h33BC	;
				14'b01101111000100: Data_out <= 16'h33B1	;
				14'b01101111000101: Data_out <= 16'h33A5	;
				14'b01101111000110: Data_out <= 16'h339A	;
				14'b01101111000111: Data_out <= 16'h338E	;
				14'b01101111001000: Data_out <= 16'h3383	;
				14'b01101111001001: Data_out <= 16'h3377	;
				14'b01101111001010: Data_out <= 16'h336C	;
				14'b01101111001011: Data_out <= 16'h3360	;
				14'b01101111001100: Data_out <= 16'h3355	;
				14'b01101111001101: Data_out <= 16'h3349	;
				14'b01101111001110: Data_out <= 16'h333E	;
				14'b01101111001111: Data_out <= 16'h3332	;
				14'b01101111010000: Data_out <= 16'h3327	;
				14'b01101111010001: Data_out <= 16'h331B	;
				14'b01101111010010: Data_out <= 16'h3310	;
				14'b01101111010011: Data_out <= 16'h3304	;
				14'b01101111010100: Data_out <= 16'h32F8	;
				14'b01101111010101: Data_out <= 16'h32ED	;
				14'b01101111010110: Data_out <= 16'h32E1	;
				14'b01101111010111: Data_out <= 16'h32D6	;
				14'b01101111011000: Data_out <= 16'h32CA	;
				14'b01101111011001: Data_out <= 16'h32BF	;
				14'b01101111011010: Data_out <= 16'h32B3	;
				14'b01101111011011: Data_out <= 16'h32A8	;
				14'b01101111011100: Data_out <= 16'h329C	;
				14'b01101111011101: Data_out <= 16'h3291	;
				14'b01101111011110: Data_out <= 16'h3285	;
				14'b01101111011111: Data_out <= 16'h327A	;
				14'b01101111100000: Data_out <= 16'h326E	;
				14'b01101111100001: Data_out <= 16'h3262	;
				14'b01101111100010: Data_out <= 16'h3257	;
				14'b01101111100011: Data_out <= 16'h324B	;
				14'b01101111100100: Data_out <= 16'h3240	;
				14'b01101111100101: Data_out <= 16'h3234	;
				14'b01101111100110: Data_out <= 16'h3229	;
				14'b01101111100111: Data_out <= 16'h321D	;
				14'b01101111101000: Data_out <= 16'h3212	;
				14'b01101111101001: Data_out <= 16'h3206	;
				14'b01101111101010: Data_out <= 16'h31FA	;
				14'b01101111101011: Data_out <= 16'h31EF	;
				14'b01101111101100: Data_out <= 16'h31E3	;
				14'b01101111101101: Data_out <= 16'h31D8	;
				14'b01101111101110: Data_out <= 16'h31CC	;
				14'b01101111101111: Data_out <= 16'h31C1	;
				14'b01101111110000: Data_out <= 16'h31B5	;
				14'b01101111110001: Data_out <= 16'h31A9	;
				14'b01101111110010: Data_out <= 16'h319E	;
				14'b01101111110011: Data_out <= 16'h3192	;
				14'b01101111110100: Data_out <= 16'h3187	;
				14'b01101111110101: Data_out <= 16'h317B	;
				14'b01101111110110: Data_out <= 16'h316F	;
				14'b01101111110111: Data_out <= 16'h3164	;
				14'b01101111111000: Data_out <= 16'h3158	;
				14'b01101111111001: Data_out <= 16'h314D	;
				14'b01101111111010: Data_out <= 16'h3141	;
				14'b01101111111011: Data_out <= 16'h3136	;
				14'b01101111111100: Data_out <= 16'h312A	;
				14'b01101111111101: Data_out <= 16'h311E	;
				14'b01101111111110: Data_out <= 16'h3113	;
				14'b01101111111111: Data_out <= 16'h3107	;
				14'b01110000000000: Data_out <= 16'h30FB	;
				14'b01110000000001: Data_out <= 16'h30F0	;
				14'b01110000000010: Data_out <= 16'h30E4	;
				14'b01110000000011: Data_out <= 16'h30D9	;
				14'b01110000000100: Data_out <= 16'h30CD	;
				14'b01110000000101: Data_out <= 16'h30C1	;
				14'b01110000000110: Data_out <= 16'h30B6	;
				14'b01110000000111: Data_out <= 16'h30AA	;
				14'b01110000001000: Data_out <= 16'h309F	;
				14'b01110000001001: Data_out <= 16'h3093	;
				14'b01110000001010: Data_out <= 16'h3087	;
				14'b01110000001011: Data_out <= 16'h307C	;
				14'b01110000001100: Data_out <= 16'h3070	;
				14'b01110000001101: Data_out <= 16'h3064	;
				14'b01110000001110: Data_out <= 16'h3059	;
				14'b01110000001111: Data_out <= 16'h304D	;
				14'b01110000010000: Data_out <= 16'h3042	;
				14'b01110000010001: Data_out <= 16'h3036	;
				14'b01110000010010: Data_out <= 16'h302A	;
				14'b01110000010011: Data_out <= 16'h301F	;
				14'b01110000010100: Data_out <= 16'h3013	;
				14'b01110000010101: Data_out <= 16'h3007	;
				14'b01110000010110: Data_out <= 16'h2FFC	;
				14'b01110000010111: Data_out <= 16'h2FF0	;
				14'b01110000011000: Data_out <= 16'h2FE4	;
				14'b01110000011001: Data_out <= 16'h2FD9	;
				14'b01110000011010: Data_out <= 16'h2FCD	;
				14'b01110000011011: Data_out <= 16'h2FC1	;
				14'b01110000011100: Data_out <= 16'h2FB6	;
				14'b01110000011101: Data_out <= 16'h2FAA	;
				14'b01110000011110: Data_out <= 16'h2F9E	;
				14'b01110000011111: Data_out <= 16'h2F93	;
				14'b01110000100000: Data_out <= 16'h2F87	;
				14'b01110000100001: Data_out <= 16'h2F7B	;
				14'b01110000100010: Data_out <= 16'h2F70	;
				14'b01110000100011: Data_out <= 16'h2F64	;
				14'b01110000100100: Data_out <= 16'h2F58	;
				14'b01110000100101: Data_out <= 16'h2F4D	;
				14'b01110000100110: Data_out <= 16'h2F41	;
				14'b01110000100111: Data_out <= 16'h2F35	;
				14'b01110000101000: Data_out <= 16'h2F2A	;
				14'b01110000101001: Data_out <= 16'h2F1E	;
				14'b01110000101010: Data_out <= 16'h2F12	;
				14'b01110000101011: Data_out <= 16'h2F07	;
				14'b01110000101100: Data_out <= 16'h2EFB	;
				14'b01110000101101: Data_out <= 16'h2EEF	;
				14'b01110000101110: Data_out <= 16'h2EE4	;
				14'b01110000101111: Data_out <= 16'h2ED8	;
				14'b01110000110000: Data_out <= 16'h2ECC	;
				14'b01110000110001: Data_out <= 16'h2EC0	;
				14'b01110000110010: Data_out <= 16'h2EB5	;
				14'b01110000110011: Data_out <= 16'h2EA9	;
				14'b01110000110100: Data_out <= 16'h2E9D	;
				14'b01110000110101: Data_out <= 16'h2E92	;
				14'b01110000110110: Data_out <= 16'h2E86	;
				14'b01110000110111: Data_out <= 16'h2E7A	;
				14'b01110000111000: Data_out <= 16'h2E6F	;
				14'b01110000111001: Data_out <= 16'h2E63	;
				14'b01110000111010: Data_out <= 16'h2E57	;
				14'b01110000111011: Data_out <= 16'h2E4B	;
				14'b01110000111100: Data_out <= 16'h2E40	;
				14'b01110000111101: Data_out <= 16'h2E34	;
				14'b01110000111110: Data_out <= 16'h2E28	;
				14'b01110000111111: Data_out <= 16'h2E1D	;
				14'b01110001000000: Data_out <= 16'h2E11	;
				14'b01110001000001: Data_out <= 16'h2E05	;
				14'b01110001000010: Data_out <= 16'h2DF9	;
				14'b01110001000011: Data_out <= 16'h2DEE	;
				14'b01110001000100: Data_out <= 16'h2DE2	;
				14'b01110001000101: Data_out <= 16'h2DD6	;
				14'b01110001000110: Data_out <= 16'h2DCA	;
				14'b01110001000111: Data_out <= 16'h2DBF	;
				14'b01110001001000: Data_out <= 16'h2DB3	;
				14'b01110001001001: Data_out <= 16'h2DA7	;
				14'b01110001001010: Data_out <= 16'h2D9B	;
				14'b01110001001011: Data_out <= 16'h2D90	;
				14'b01110001001100: Data_out <= 16'h2D84	;
				14'b01110001001101: Data_out <= 16'h2D78	;
				14'b01110001001110: Data_out <= 16'h2D6C	;
				14'b01110001001111: Data_out <= 16'h2D61	;
				14'b01110001010000: Data_out <= 16'h2D55	;
				14'b01110001010001: Data_out <= 16'h2D49	;
				14'b01110001010010: Data_out <= 16'h2D3D	;
				14'b01110001010011: Data_out <= 16'h2D32	;
				14'b01110001010100: Data_out <= 16'h2D26	;
				14'b01110001010101: Data_out <= 16'h2D1A	;
				14'b01110001010110: Data_out <= 16'h2D0E	;
				14'b01110001010111: Data_out <= 16'h2D03	;
				14'b01110001011000: Data_out <= 16'h2CF7	;
				14'b01110001011001: Data_out <= 16'h2CEB	;
				14'b01110001011010: Data_out <= 16'h2CDF	;
				14'b01110001011011: Data_out <= 16'h2CD4	;
				14'b01110001011100: Data_out <= 16'h2CC8	;
				14'b01110001011101: Data_out <= 16'h2CBC	;
				14'b01110001011110: Data_out <= 16'h2CB0	;
				14'b01110001011111: Data_out <= 16'h2CA5	;
				14'b01110001100000: Data_out <= 16'h2C99	;
				14'b01110001100001: Data_out <= 16'h2C8D	;
				14'b01110001100010: Data_out <= 16'h2C81	;
				14'b01110001100011: Data_out <= 16'h2C75	;
				14'b01110001100100: Data_out <= 16'h2C6A	;
				14'b01110001100101: Data_out <= 16'h2C5E	;
				14'b01110001100110: Data_out <= 16'h2C52	;
				14'b01110001100111: Data_out <= 16'h2C46	;
				14'b01110001101000: Data_out <= 16'h2C3A	;
				14'b01110001101001: Data_out <= 16'h2C2F	;
				14'b01110001101010: Data_out <= 16'h2C23	;
				14'b01110001101011: Data_out <= 16'h2C17	;
				14'b01110001101100: Data_out <= 16'h2C0B	;
				14'b01110001101101: Data_out <= 16'h2BFF	;
				14'b01110001101110: Data_out <= 16'h2BF4	;
				14'b01110001101111: Data_out <= 16'h2BE8	;
				14'b01110001110000: Data_out <= 16'h2BDC	;
				14'b01110001110001: Data_out <= 16'h2BD0	;
				14'b01110001110010: Data_out <= 16'h2BC4	;
				14'b01110001110011: Data_out <= 16'h2BB9	;
				14'b01110001110100: Data_out <= 16'h2BAD	;
				14'b01110001110101: Data_out <= 16'h2BA1	;
				14'b01110001110110: Data_out <= 16'h2B95	;
				14'b01110001110111: Data_out <= 16'h2B89	;
				14'b01110001111000: Data_out <= 16'h2B7E	;
				14'b01110001111001: Data_out <= 16'h2B72	;
				14'b01110001111010: Data_out <= 16'h2B66	;
				14'b01110001111011: Data_out <= 16'h2B5A	;
				14'b01110001111100: Data_out <= 16'h2B4E	;
				14'b01110001111101: Data_out <= 16'h2B42	;
				14'b01110001111110: Data_out <= 16'h2B37	;
				14'b01110001111111: Data_out <= 16'h2B2B	;
				14'b01110010000000: Data_out <= 16'h2B1F	;
				14'b01110010000001: Data_out <= 16'h2B13	;
				14'b01110010000010: Data_out <= 16'h2B07	;
				14'b01110010000011: Data_out <= 16'h2AFB	;
				14'b01110010000100: Data_out <= 16'h2AF0	;
				14'b01110010000101: Data_out <= 16'h2AE4	;
				14'b01110010000110: Data_out <= 16'h2AD8	;
				14'b01110010000111: Data_out <= 16'h2ACC	;
				14'b01110010001000: Data_out <= 16'h2AC0	;
				14'b01110010001001: Data_out <= 16'h2AB4	;
				14'b01110010001010: Data_out <= 16'h2AA9	;
				14'b01110010001011: Data_out <= 16'h2A9D	;
				14'b01110010001100: Data_out <= 16'h2A91	;
				14'b01110010001101: Data_out <= 16'h2A85	;
				14'b01110010001110: Data_out <= 16'h2A79	;
				14'b01110010001111: Data_out <= 16'h2A6D	;
				14'b01110010010000: Data_out <= 16'h2A61	;
				14'b01110010010001: Data_out <= 16'h2A56	;
				14'b01110010010010: Data_out <= 16'h2A4A	;
				14'b01110010010011: Data_out <= 16'h2A3E	;
				14'b01110010010100: Data_out <= 16'h2A32	;
				14'b01110010010101: Data_out <= 16'h2A26	;
				14'b01110010010110: Data_out <= 16'h2A1A	;
				14'b01110010010111: Data_out <= 16'h2A0E	;
				14'b01110010011000: Data_out <= 16'h2A03	;
				14'b01110010011001: Data_out <= 16'h29F7	;
				14'b01110010011010: Data_out <= 16'h29EB	;
				14'b01110010011011: Data_out <= 16'h29DF	;
				14'b01110010011100: Data_out <= 16'h29D3	;
				14'b01110010011101: Data_out <= 16'h29C7	;
				14'b01110010011110: Data_out <= 16'h29BB	;
				14'b01110010011111: Data_out <= 16'h29AF	;
				14'b01110010100000: Data_out <= 16'h29A4	;
				14'b01110010100001: Data_out <= 16'h2998	;
				14'b01110010100010: Data_out <= 16'h298C	;
				14'b01110010100011: Data_out <= 16'h2980	;
				14'b01110010100100: Data_out <= 16'h2974	;
				14'b01110010100101: Data_out <= 16'h2968	;
				14'b01110010100110: Data_out <= 16'h295C	;
				14'b01110010100111: Data_out <= 16'h2950	;
				14'b01110010101000: Data_out <= 16'h2944	;
				14'b01110010101001: Data_out <= 16'h2939	;
				14'b01110010101010: Data_out <= 16'h292D	;
				14'b01110010101011: Data_out <= 16'h2921	;
				14'b01110010101100: Data_out <= 16'h2915	;
				14'b01110010101101: Data_out <= 16'h2909	;
				14'b01110010101110: Data_out <= 16'h28FD	;
				14'b01110010101111: Data_out <= 16'h28F1	;
				14'b01110010110000: Data_out <= 16'h28E5	;
				14'b01110010110001: Data_out <= 16'h28D9	;
				14'b01110010110010: Data_out <= 16'h28CD	;
				14'b01110010110011: Data_out <= 16'h28C1	;
				14'b01110010110100: Data_out <= 16'h28B6	;
				14'b01110010110101: Data_out <= 16'h28AA	;
				14'b01110010110110: Data_out <= 16'h289E	;
				14'b01110010110111: Data_out <= 16'h2892	;
				14'b01110010111000: Data_out <= 16'h2886	;
				14'b01110010111001: Data_out <= 16'h287A	;
				14'b01110010111010: Data_out <= 16'h286E	;
				14'b01110010111011: Data_out <= 16'h2862	;
				14'b01110010111100: Data_out <= 16'h2856	;
				14'b01110010111101: Data_out <= 16'h284A	;
				14'b01110010111110: Data_out <= 16'h283E	;
				14'b01110010111111: Data_out <= 16'h2832	;
				14'b01110011000000: Data_out <= 16'h2827	;
				14'b01110011000001: Data_out <= 16'h281B	;
				14'b01110011000010: Data_out <= 16'h280F	;
				14'b01110011000011: Data_out <= 16'h2803	;
				14'b01110011000100: Data_out <= 16'h27F7	;
				14'b01110011000101: Data_out <= 16'h27EB	;
				14'b01110011000110: Data_out <= 16'h27DF	;
				14'b01110011000111: Data_out <= 16'h27D3	;
				14'b01110011001000: Data_out <= 16'h27C7	;
				14'b01110011001001: Data_out <= 16'h27BB	;
				14'b01110011001010: Data_out <= 16'h27AF	;
				14'b01110011001011: Data_out <= 16'h27A3	;
				14'b01110011001100: Data_out <= 16'h2797	;
				14'b01110011001101: Data_out <= 16'h278B	;
				14'b01110011001110: Data_out <= 16'h277F	;
				14'b01110011001111: Data_out <= 16'h2773	;
				14'b01110011010000: Data_out <= 16'h2767	;
				14'b01110011010001: Data_out <= 16'h275B	;
				14'b01110011010010: Data_out <= 16'h274F	;
				14'b01110011010011: Data_out <= 16'h2744	;
				14'b01110011010100: Data_out <= 16'h2738	;
				14'b01110011010101: Data_out <= 16'h272C	;
				14'b01110011010110: Data_out <= 16'h2720	;
				14'b01110011010111: Data_out <= 16'h2714	;
				14'b01110011011000: Data_out <= 16'h2708	;
				14'b01110011011001: Data_out <= 16'h26FC	;
				14'b01110011011010: Data_out <= 16'h26F0	;
				14'b01110011011011: Data_out <= 16'h26E4	;
				14'b01110011011100: Data_out <= 16'h26D8	;
				14'b01110011011101: Data_out <= 16'h26CC	;
				14'b01110011011110: Data_out <= 16'h26C0	;
				14'b01110011011111: Data_out <= 16'h26B4	;
				14'b01110011100000: Data_out <= 16'h26A8	;
				14'b01110011100001: Data_out <= 16'h269C	;
				14'b01110011100010: Data_out <= 16'h2690	;
				14'b01110011100011: Data_out <= 16'h2684	;
				14'b01110011100100: Data_out <= 16'h2678	;
				14'b01110011100101: Data_out <= 16'h266C	;
				14'b01110011100110: Data_out <= 16'h2660	;
				14'b01110011100111: Data_out <= 16'h2654	;
				14'b01110011101000: Data_out <= 16'h2648	;
				14'b01110011101001: Data_out <= 16'h263C	;
				14'b01110011101010: Data_out <= 16'h2630	;
				14'b01110011101011: Data_out <= 16'h2624	;
				14'b01110011101100: Data_out <= 16'h2618	;
				14'b01110011101101: Data_out <= 16'h260C	;
				14'b01110011101110: Data_out <= 16'h2600	;
				14'b01110011101111: Data_out <= 16'h25F4	;
				14'b01110011110000: Data_out <= 16'h25E8	;
				14'b01110011110001: Data_out <= 16'h25DC	;
				14'b01110011110010: Data_out <= 16'h25D0	;
				14'b01110011110011: Data_out <= 16'h25C4	;
				14'b01110011110100: Data_out <= 16'h25B8	;
				14'b01110011110101: Data_out <= 16'h25AC	;
				14'b01110011110110: Data_out <= 16'h25A0	;
				14'b01110011110111: Data_out <= 16'h2594	;
				14'b01110011111000: Data_out <= 16'h2588	;
				14'b01110011111001: Data_out <= 16'h257C	;
				14'b01110011111010: Data_out <= 16'h2570	;
				14'b01110011111011: Data_out <= 16'h2564	;
				14'b01110011111100: Data_out <= 16'h2558	;
				14'b01110011111101: Data_out <= 16'h254C	;
				14'b01110011111110: Data_out <= 16'h2540	;
				14'b01110011111111: Data_out <= 16'h2534	;
				14'b01110100000000: Data_out <= 16'h2528	;
				14'b01110100000001: Data_out <= 16'h251C	;
				14'b01110100000010: Data_out <= 16'h2510	;
				14'b01110100000011: Data_out <= 16'h2504	;
				14'b01110100000100: Data_out <= 16'h24F8	;
				14'b01110100000101: Data_out <= 16'h24EC	;
				14'b01110100000110: Data_out <= 16'h24E0	;
				14'b01110100000111: Data_out <= 16'h24D4	;
				14'b01110100001000: Data_out <= 16'h24C8	;
				14'b01110100001001: Data_out <= 16'h24BC	;
				14'b01110100001010: Data_out <= 16'h24B0	;
				14'b01110100001011: Data_out <= 16'h24A3	;
				14'b01110100001100: Data_out <= 16'h2497	;
				14'b01110100001101: Data_out <= 16'h248B	;
				14'b01110100001110: Data_out <= 16'h247F	;
				14'b01110100001111: Data_out <= 16'h2473	;
				14'b01110100010000: Data_out <= 16'h2467	;
				14'b01110100010001: Data_out <= 16'h245B	;
				14'b01110100010010: Data_out <= 16'h244F	;
				14'b01110100010011: Data_out <= 16'h2443	;
				14'b01110100010100: Data_out <= 16'h2437	;
				14'b01110100010101: Data_out <= 16'h242B	;
				14'b01110100010110: Data_out <= 16'h241F	;
				14'b01110100010111: Data_out <= 16'h2413	;
				14'b01110100011000: Data_out <= 16'h2407	;
				14'b01110100011001: Data_out <= 16'h23FB	;
				14'b01110100011010: Data_out <= 16'h23EF	;
				14'b01110100011011: Data_out <= 16'h23E3	;
				14'b01110100011100: Data_out <= 16'h23D7	;
				14'b01110100011101: Data_out <= 16'h23CB	;
				14'b01110100011110: Data_out <= 16'h23BE	;
				14'b01110100011111: Data_out <= 16'h23B2	;
				14'b01110100100000: Data_out <= 16'h23A6	;
				14'b01110100100001: Data_out <= 16'h239A	;
				14'b01110100100010: Data_out <= 16'h238E	;
				14'b01110100100011: Data_out <= 16'h2382	;
				14'b01110100100100: Data_out <= 16'h2376	;
				14'b01110100100101: Data_out <= 16'h236A	;
				14'b01110100100110: Data_out <= 16'h235E	;
				14'b01110100100111: Data_out <= 16'h2352	;
				14'b01110100101000: Data_out <= 16'h2346	;
				14'b01110100101001: Data_out <= 16'h233A	;
				14'b01110100101010: Data_out <= 16'h232E	;
				14'b01110100101011: Data_out <= 16'h2322	;
				14'b01110100101100: Data_out <= 16'h2315	;
				14'b01110100101101: Data_out <= 16'h2309	;
				14'b01110100101110: Data_out <= 16'h22FD	;
				14'b01110100101111: Data_out <= 16'h22F1	;
				14'b01110100110000: Data_out <= 16'h22E5	;
				14'b01110100110001: Data_out <= 16'h22D9	;
				14'b01110100110010: Data_out <= 16'h22CD	;
				14'b01110100110011: Data_out <= 16'h22C1	;
				14'b01110100110100: Data_out <= 16'h22B5	;
				14'b01110100110101: Data_out <= 16'h22A9	;
				14'b01110100110110: Data_out <= 16'h229D	;
				14'b01110100110111: Data_out <= 16'h2290	;
				14'b01110100111000: Data_out <= 16'h2284	;
				14'b01110100111001: Data_out <= 16'h2278	;
				14'b01110100111010: Data_out <= 16'h226C	;
				14'b01110100111011: Data_out <= 16'h2260	;
				14'b01110100111100: Data_out <= 16'h2254	;
				14'b01110100111101: Data_out <= 16'h2248	;
				14'b01110100111110: Data_out <= 16'h223C	;
				14'b01110100111111: Data_out <= 16'h2230	;
				14'b01110101000000: Data_out <= 16'h2223	;
				14'b01110101000001: Data_out <= 16'h2217	;
				14'b01110101000010: Data_out <= 16'h220B	;
				14'b01110101000011: Data_out <= 16'h21FF	;
				14'b01110101000100: Data_out <= 16'h21F3	;
				14'b01110101000101: Data_out <= 16'h21E7	;
				14'b01110101000110: Data_out <= 16'h21DB	;
				14'b01110101000111: Data_out <= 16'h21CF	;
				14'b01110101001000: Data_out <= 16'h21C3	;
				14'b01110101001001: Data_out <= 16'h21B6	;
				14'b01110101001010: Data_out <= 16'h21AA	;
				14'b01110101001011: Data_out <= 16'h219E	;
				14'b01110101001100: Data_out <= 16'h2192	;
				14'b01110101001101: Data_out <= 16'h2186	;
				14'b01110101001110: Data_out <= 16'h217A	;
				14'b01110101001111: Data_out <= 16'h216E	;
				14'b01110101010000: Data_out <= 16'h2162	;
				14'b01110101010001: Data_out <= 16'h2155	;
				14'b01110101010010: Data_out <= 16'h2149	;
				14'b01110101010011: Data_out <= 16'h213D	;
				14'b01110101010100: Data_out <= 16'h2131	;
				14'b01110101010101: Data_out <= 16'h2125	;
				14'b01110101010110: Data_out <= 16'h2119	;
				14'b01110101010111: Data_out <= 16'h210D	;
				14'b01110101011000: Data_out <= 16'h2100	;
				14'b01110101011001: Data_out <= 16'h20F4	;
				14'b01110101011010: Data_out <= 16'h20E8	;
				14'b01110101011011: Data_out <= 16'h20DC	;
				14'b01110101011100: Data_out <= 16'h20D0	;
				14'b01110101011101: Data_out <= 16'h20C4	;
				14'b01110101011110: Data_out <= 16'h20B8	;
				14'b01110101011111: Data_out <= 16'h20AB	;
				14'b01110101100000: Data_out <= 16'h209F	;
				14'b01110101100001: Data_out <= 16'h2093	;
				14'b01110101100010: Data_out <= 16'h2087	;
				14'b01110101100011: Data_out <= 16'h207B	;
				14'b01110101100100: Data_out <= 16'h206F	;
				14'b01110101100101: Data_out <= 16'h2063	;
				14'b01110101100110: Data_out <= 16'h2056	;
				14'b01110101100111: Data_out <= 16'h204A	;
				14'b01110101101000: Data_out <= 16'h203E	;
				14'b01110101101001: Data_out <= 16'h2032	;
				14'b01110101101010: Data_out <= 16'h2026	;
				14'b01110101101011: Data_out <= 16'h201A	;
				14'b01110101101100: Data_out <= 16'h200D	;
				14'b01110101101101: Data_out <= 16'h2001	;
				14'b01110101101110: Data_out <= 16'h1FF5	;
				14'b01110101101111: Data_out <= 16'h1FE9	;
				14'b01110101110000: Data_out <= 16'h1FDD	;
				14'b01110101110001: Data_out <= 16'h1FD1	;
				14'b01110101110010: Data_out <= 16'h1FC4	;
				14'b01110101110011: Data_out <= 16'h1FB8	;
				14'b01110101110100: Data_out <= 16'h1FAC	;
				14'b01110101110101: Data_out <= 16'h1FA0	;
				14'b01110101110110: Data_out <= 16'h1F94	;
				14'b01110101110111: Data_out <= 16'h1F87	;
				14'b01110101111000: Data_out <= 16'h1F7B	;
				14'b01110101111001: Data_out <= 16'h1F6F	;
				14'b01110101111010: Data_out <= 16'h1F63	;
				14'b01110101111011: Data_out <= 16'h1F57	;
				14'b01110101111100: Data_out <= 16'h1F4B	;
				14'b01110101111101: Data_out <= 16'h1F3E	;
				14'b01110101111110: Data_out <= 16'h1F32	;
				14'b01110101111111: Data_out <= 16'h1F26	;
				14'b01110110000000: Data_out <= 16'h1F1A	;
				14'b01110110000001: Data_out <= 16'h1F0E	;
				14'b01110110000010: Data_out <= 16'h1F01	;
				14'b01110110000011: Data_out <= 16'h1EF5	;
				14'b01110110000100: Data_out <= 16'h1EE9	;
				14'b01110110000101: Data_out <= 16'h1EDD	;
				14'b01110110000110: Data_out <= 16'h1ED1	;
				14'b01110110000111: Data_out <= 16'h1EC4	;
				14'b01110110001000: Data_out <= 16'h1EB8	;
				14'b01110110001001: Data_out <= 16'h1EAC	;
				14'b01110110001010: Data_out <= 16'h1EA0	;
				14'b01110110001011: Data_out <= 16'h1E94	;
				14'b01110110001100: Data_out <= 16'h1E87	;
				14'b01110110001101: Data_out <= 16'h1E7B	;
				14'b01110110001110: Data_out <= 16'h1E6F	;
				14'b01110110001111: Data_out <= 16'h1E63	;
				14'b01110110010000: Data_out <= 16'h1E57	;
				14'b01110110010001: Data_out <= 16'h1E4A	;
				14'b01110110010010: Data_out <= 16'h1E3E	;
				14'b01110110010011: Data_out <= 16'h1E32	;
				14'b01110110010100: Data_out <= 16'h1E26	;
				14'b01110110010101: Data_out <= 16'h1E1A	;
				14'b01110110010110: Data_out <= 16'h1E0D	;
				14'b01110110010111: Data_out <= 16'h1E01	;
				14'b01110110011000: Data_out <= 16'h1DF5	;
				14'b01110110011001: Data_out <= 16'h1DE9	;
				14'b01110110011010: Data_out <= 16'h1DDD	;
				14'b01110110011011: Data_out <= 16'h1DD0	;
				14'b01110110011100: Data_out <= 16'h1DC4	;
				14'b01110110011101: Data_out <= 16'h1DB8	;
				14'b01110110011110: Data_out <= 16'h1DAC	;
				14'b01110110011111: Data_out <= 16'h1D9F	;
				14'b01110110100000: Data_out <= 16'h1D93	;
				14'b01110110100001: Data_out <= 16'h1D87	;
				14'b01110110100010: Data_out <= 16'h1D7B	;
				14'b01110110100011: Data_out <= 16'h1D6E	;
				14'b01110110100100: Data_out <= 16'h1D62	;
				14'b01110110100101: Data_out <= 16'h1D56	;
				14'b01110110100110: Data_out <= 16'h1D4A	;
				14'b01110110100111: Data_out <= 16'h1D3E	;
				14'b01110110101000: Data_out <= 16'h1D31	;
				14'b01110110101001: Data_out <= 16'h1D25	;
				14'b01110110101010: Data_out <= 16'h1D19	;
				14'b01110110101011: Data_out <= 16'h1D0D	;
				14'b01110110101100: Data_out <= 16'h1D00	;
				14'b01110110101101: Data_out <= 16'h1CF4	;
				14'b01110110101110: Data_out <= 16'h1CE8	;
				14'b01110110101111: Data_out <= 16'h1CDC	;
				14'b01110110110000: Data_out <= 16'h1CCF	;
				14'b01110110110001: Data_out <= 16'h1CC3	;
				14'b01110110110010: Data_out <= 16'h1CB7	;
				14'b01110110110011: Data_out <= 16'h1CAB	;
				14'b01110110110100: Data_out <= 16'h1C9E	;
				14'b01110110110101: Data_out <= 16'h1C92	;
				14'b01110110110110: Data_out <= 16'h1C86	;
				14'b01110110110111: Data_out <= 16'h1C7A	;
				14'b01110110111000: Data_out <= 16'h1C6D	;
				14'b01110110111001: Data_out <= 16'h1C61	;
				14'b01110110111010: Data_out <= 16'h1C55	;
				14'b01110110111011: Data_out <= 16'h1C49	;
				14'b01110110111100: Data_out <= 16'h1C3C	;
				14'b01110110111101: Data_out <= 16'h1C30	;
				14'b01110110111110: Data_out <= 16'h1C24	;
				14'b01110110111111: Data_out <= 16'h1C18	;
				14'b01110111000000: Data_out <= 16'h1C0B	;
				14'b01110111000001: Data_out <= 16'h1BFF	;
				14'b01110111000010: Data_out <= 16'h1BF3	;
				14'b01110111000011: Data_out <= 16'h1BE7	;
				14'b01110111000100: Data_out <= 16'h1BDA	;
				14'b01110111000101: Data_out <= 16'h1BCE	;
				14'b01110111000110: Data_out <= 16'h1BC2	;
				14'b01110111000111: Data_out <= 16'h1BB6	;
				14'b01110111001000: Data_out <= 16'h1BA9	;
				14'b01110111001001: Data_out <= 16'h1B9D	;
				14'b01110111001010: Data_out <= 16'h1B91	;
				14'b01110111001011: Data_out <= 16'h1B84	;
				14'b01110111001100: Data_out <= 16'h1B78	;
				14'b01110111001101: Data_out <= 16'h1B6C	;
				14'b01110111001110: Data_out <= 16'h1B60	;
				14'b01110111001111: Data_out <= 16'h1B53	;
				14'b01110111010000: Data_out <= 16'h1B47	;
				14'b01110111010001: Data_out <= 16'h1B3B	;
				14'b01110111010010: Data_out <= 16'h1B2F	;
				14'b01110111010011: Data_out <= 16'h1B22	;
				14'b01110111010100: Data_out <= 16'h1B16	;
				14'b01110111010101: Data_out <= 16'h1B0A	;
				14'b01110111010110: Data_out <= 16'h1AFD	;
				14'b01110111010111: Data_out <= 16'h1AF1	;
				14'b01110111011000: Data_out <= 16'h1AE5	;
				14'b01110111011001: Data_out <= 16'h1AD9	;
				14'b01110111011010: Data_out <= 16'h1ACC	;
				14'b01110111011011: Data_out <= 16'h1AC0	;
				14'b01110111011100: Data_out <= 16'h1AB4	;
				14'b01110111011101: Data_out <= 16'h1AA7	;
				14'b01110111011110: Data_out <= 16'h1A9B	;
				14'b01110111011111: Data_out <= 16'h1A8F	;
				14'b01110111100000: Data_out <= 16'h1A83	;
				14'b01110111100001: Data_out <= 16'h1A76	;
				14'b01110111100010: Data_out <= 16'h1A6A	;
				14'b01110111100011: Data_out <= 16'h1A5E	;
				14'b01110111100100: Data_out <= 16'h1A51	;
				14'b01110111100101: Data_out <= 16'h1A45	;
				14'b01110111100110: Data_out <= 16'h1A39	;
				14'b01110111100111: Data_out <= 16'h1A2C	;
				14'b01110111101000: Data_out <= 16'h1A20	;
				14'b01110111101001: Data_out <= 16'h1A14	;
				14'b01110111101010: Data_out <= 16'h1A08	;
				14'b01110111101011: Data_out <= 16'h19FB	;
				14'b01110111101100: Data_out <= 16'h19EF	;
				14'b01110111101101: Data_out <= 16'h19E3	;
				14'b01110111101110: Data_out <= 16'h19D6	;
				14'b01110111101111: Data_out <= 16'h19CA	;
				14'b01110111110000: Data_out <= 16'h19BE	;
				14'b01110111110001: Data_out <= 16'h19B1	;
				14'b01110111110010: Data_out <= 16'h19A5	;
				14'b01110111110011: Data_out <= 16'h1999	;
				14'b01110111110100: Data_out <= 16'h198C	;
				14'b01110111110101: Data_out <= 16'h1980	;
				14'b01110111110110: Data_out <= 16'h1974	;
				14'b01110111110111: Data_out <= 16'h1968	;
				14'b01110111111000: Data_out <= 16'h195B	;
				14'b01110111111001: Data_out <= 16'h194F	;
				14'b01110111111010: Data_out <= 16'h1943	;
				14'b01110111111011: Data_out <= 16'h1936	;
				14'b01110111111100: Data_out <= 16'h192A	;
				14'b01110111111101: Data_out <= 16'h191E	;
				14'b01110111111110: Data_out <= 16'h1911	;
				14'b01110111111111: Data_out <= 16'h1905	;
				14'b01111000000000: Data_out <= 16'h18F9	;
				14'b01111000000001: Data_out <= 16'h18EC	;
				14'b01111000000010: Data_out <= 16'h18E0	;
				14'b01111000000011: Data_out <= 16'h18D4	;
				14'b01111000000100: Data_out <= 16'h18C7	;
				14'b01111000000101: Data_out <= 16'h18BB	;
				14'b01111000000110: Data_out <= 16'h18AF	;
				14'b01111000000111: Data_out <= 16'h18A2	;
				14'b01111000001000: Data_out <= 16'h1896	;
				14'b01111000001001: Data_out <= 16'h188A	;
				14'b01111000001010: Data_out <= 16'h187D	;
				14'b01111000001011: Data_out <= 16'h1871	;
				14'b01111000001100: Data_out <= 16'h1865	;
				14'b01111000001101: Data_out <= 16'h1858	;
				14'b01111000001110: Data_out <= 16'h184C	;
				14'b01111000001111: Data_out <= 16'h1840	;
				14'b01111000010000: Data_out <= 16'h1833	;
				14'b01111000010001: Data_out <= 16'h1827	;
				14'b01111000010010: Data_out <= 16'h181B	;
				14'b01111000010011: Data_out <= 16'h180E	;
				14'b01111000010100: Data_out <= 16'h1802	;
				14'b01111000010101: Data_out <= 16'h17F6	;
				14'b01111000010110: Data_out <= 16'h17E9	;
				14'b01111000010111: Data_out <= 16'h17DD	;
				14'b01111000011000: Data_out <= 16'h17D1	;
				14'b01111000011001: Data_out <= 16'h17C4	;
				14'b01111000011010: Data_out <= 16'h17B8	;
				14'b01111000011011: Data_out <= 16'h17AC	;
				14'b01111000011100: Data_out <= 16'h179F	;
				14'b01111000011101: Data_out <= 16'h1793	;
				14'b01111000011110: Data_out <= 16'h1786	;
				14'b01111000011111: Data_out <= 16'h177A	;
				14'b01111000100000: Data_out <= 16'h176E	;
				14'b01111000100001: Data_out <= 16'h1761	;
				14'b01111000100010: Data_out <= 16'h1755	;
				14'b01111000100011: Data_out <= 16'h1749	;
				14'b01111000100100: Data_out <= 16'h173C	;
				14'b01111000100101: Data_out <= 16'h1730	;
				14'b01111000100110: Data_out <= 16'h1724	;
				14'b01111000100111: Data_out <= 16'h1717	;
				14'b01111000101000: Data_out <= 16'h170B	;
				14'b01111000101001: Data_out <= 16'h16FF	;
				14'b01111000101010: Data_out <= 16'h16F2	;
				14'b01111000101011: Data_out <= 16'h16E6	;
				14'b01111000101100: Data_out <= 16'h16D9	;
				14'b01111000101101: Data_out <= 16'h16CD	;
				14'b01111000101110: Data_out <= 16'h16C1	;
				14'b01111000101111: Data_out <= 16'h16B4	;
				14'b01111000110000: Data_out <= 16'h16A8	;
				14'b01111000110001: Data_out <= 16'h169C	;
				14'b01111000110010: Data_out <= 16'h168F	;
				14'b01111000110011: Data_out <= 16'h1683	;
				14'b01111000110100: Data_out <= 16'h1677	;
				14'b01111000110101: Data_out <= 16'h166A	;
				14'b01111000110110: Data_out <= 16'h165E	;
				14'b01111000110111: Data_out <= 16'h1651	;
				14'b01111000111000: Data_out <= 16'h1645	;
				14'b01111000111001: Data_out <= 16'h1639	;
				14'b01111000111010: Data_out <= 16'h162C	;
				14'b01111000111011: Data_out <= 16'h1620	;
				14'b01111000111100: Data_out <= 16'h1614	;
				14'b01111000111101: Data_out <= 16'h1607	;
				14'b01111000111110: Data_out <= 16'h15FB	;
				14'b01111000111111: Data_out <= 16'h15EE	;
				14'b01111001000000: Data_out <= 16'h15E2	;
				14'b01111001000001: Data_out <= 16'h15D6	;
				14'b01111001000010: Data_out <= 16'h15C9	;
				14'b01111001000011: Data_out <= 16'h15BD	;
				14'b01111001000100: Data_out <= 16'h15B0	;
				14'b01111001000101: Data_out <= 16'h15A4	;
				14'b01111001000110: Data_out <= 16'h1598	;
				14'b01111001000111: Data_out <= 16'h158B	;
				14'b01111001001000: Data_out <= 16'h157F	;
				14'b01111001001001: Data_out <= 16'h1573	;
				14'b01111001001010: Data_out <= 16'h1566	;
				14'b01111001001011: Data_out <= 16'h155A	;
				14'b01111001001100: Data_out <= 16'h154D	;
				14'b01111001001101: Data_out <= 16'h1541	;
				14'b01111001001110: Data_out <= 16'h1535	;
				14'b01111001001111: Data_out <= 16'h1528	;
				14'b01111001010000: Data_out <= 16'h151C	;
				14'b01111001010001: Data_out <= 16'h150F	;
				14'b01111001010010: Data_out <= 16'h1503	;
				14'b01111001010011: Data_out <= 16'h14F7	;
				14'b01111001010100: Data_out <= 16'h14EA	;
				14'b01111001010101: Data_out <= 16'h14DE	;
				14'b01111001010110: Data_out <= 16'h14D1	;
				14'b01111001010111: Data_out <= 16'h14C5	;
				14'b01111001011000: Data_out <= 16'h14B9	;
				14'b01111001011001: Data_out <= 16'h14AC	;
				14'b01111001011010: Data_out <= 16'h14A0	;
				14'b01111001011011: Data_out <= 16'h1493	;
				14'b01111001011100: Data_out <= 16'h1487	;
				14'b01111001011101: Data_out <= 16'h147B	;
				14'b01111001011110: Data_out <= 16'h146E	;
				14'b01111001011111: Data_out <= 16'h1462	;
				14'b01111001100000: Data_out <= 16'h1455	;
				14'b01111001100001: Data_out <= 16'h1449	;
				14'b01111001100010: Data_out <= 16'h143D	;
				14'b01111001100011: Data_out <= 16'h1430	;
				14'b01111001100100: Data_out <= 16'h1424	;
				14'b01111001100101: Data_out <= 16'h1417	;
				14'b01111001100110: Data_out <= 16'h140B	;
				14'b01111001100111: Data_out <= 16'h13FF	;
				14'b01111001101000: Data_out <= 16'h13F2	;
				14'b01111001101001: Data_out <= 16'h13E6	;
				14'b01111001101010: Data_out <= 16'h13D9	;
				14'b01111001101011: Data_out <= 16'h13CD	;
				14'b01111001101100: Data_out <= 16'h13C0	;
				14'b01111001101101: Data_out <= 16'h13B4	;
				14'b01111001101110: Data_out <= 16'h13A8	;
				14'b01111001101111: Data_out <= 16'h139B	;
				14'b01111001110000: Data_out <= 16'h138F	;
				14'b01111001110001: Data_out <= 16'h1382	;
				14'b01111001110010: Data_out <= 16'h1376	;
				14'b01111001110011: Data_out <= 16'h136A	;
				14'b01111001110100: Data_out <= 16'h135D	;
				14'b01111001110101: Data_out <= 16'h1351	;
				14'b01111001110110: Data_out <= 16'h1344	;
				14'b01111001110111: Data_out <= 16'h1338	;
				14'b01111001111000: Data_out <= 16'h132B	;
				14'b01111001111001: Data_out <= 16'h131F	;
				14'b01111001111010: Data_out <= 16'h1313	;
				14'b01111001111011: Data_out <= 16'h1306	;
				14'b01111001111100: Data_out <= 16'h12FA	;
				14'b01111001111101: Data_out <= 16'h12ED	;
				14'b01111001111110: Data_out <= 16'h12E1	;
				14'b01111001111111: Data_out <= 16'h12D4	;
				14'b01111010000000: Data_out <= 16'h12C8	;
				14'b01111010000001: Data_out <= 16'h12BC	;
				14'b01111010000010: Data_out <= 16'h12AF	;
				14'b01111010000011: Data_out <= 16'h12A3	;
				14'b01111010000100: Data_out <= 16'h1296	;
				14'b01111010000101: Data_out <= 16'h128A	;
				14'b01111010000110: Data_out <= 16'h127D	;
				14'b01111010000111: Data_out <= 16'h1271	;
				14'b01111010001000: Data_out <= 16'h1265	;
				14'b01111010001001: Data_out <= 16'h1258	;
				14'b01111010001010: Data_out <= 16'h124C	;
				14'b01111010001011: Data_out <= 16'h123F	;
				14'b01111010001100: Data_out <= 16'h1233	;
				14'b01111010001101: Data_out <= 16'h1226	;
				14'b01111010001110: Data_out <= 16'h121A	;
				14'b01111010001111: Data_out <= 16'h120D	;
				14'b01111010010000: Data_out <= 16'h1201	;
				14'b01111010010001: Data_out <= 16'h11F5	;
				14'b01111010010010: Data_out <= 16'h11E8	;
				14'b01111010010011: Data_out <= 16'h11DC	;
				14'b01111010010100: Data_out <= 16'h11CF	;
				14'b01111010010101: Data_out <= 16'h11C3	;
				14'b01111010010110: Data_out <= 16'h11B6	;
				14'b01111010010111: Data_out <= 16'h11AA	;
				14'b01111010011000: Data_out <= 16'h119D	;
				14'b01111010011001: Data_out <= 16'h1191	;
				14'b01111010011010: Data_out <= 16'h1185	;
				14'b01111010011011: Data_out <= 16'h1178	;
				14'b01111010011100: Data_out <= 16'h116C	;
				14'b01111010011101: Data_out <= 16'h115F	;
				14'b01111010011110: Data_out <= 16'h1153	;
				14'b01111010011111: Data_out <= 16'h1146	;
				14'b01111010100000: Data_out <= 16'h113A	;
				14'b01111010100001: Data_out <= 16'h112D	;
				14'b01111010100010: Data_out <= 16'h1121	;
				14'b01111010100011: Data_out <= 16'h1115	;
				14'b01111010100100: Data_out <= 16'h1108	;
				14'b01111010100101: Data_out <= 16'h10FC	;
				14'b01111010100110: Data_out <= 16'h10EF	;
				14'b01111010100111: Data_out <= 16'h10E3	;
				14'b01111010101000: Data_out <= 16'h10D6	;
				14'b01111010101001: Data_out <= 16'h10CA	;
				14'b01111010101010: Data_out <= 16'h10BD	;
				14'b01111010101011: Data_out <= 16'h10B1	;
				14'b01111010101100: Data_out <= 16'h10A4	;
				14'b01111010101101: Data_out <= 16'h1098	;
				14'b01111010101110: Data_out <= 16'h108C	;
				14'b01111010101111: Data_out <= 16'h107F	;
				14'b01111010110000: Data_out <= 16'h1073	;
				14'b01111010110001: Data_out <= 16'h1066	;
				14'b01111010110010: Data_out <= 16'h105A	;
				14'b01111010110011: Data_out <= 16'h104D	;
				14'b01111010110100: Data_out <= 16'h1041	;
				14'b01111010110101: Data_out <= 16'h1034	;
				14'b01111010110110: Data_out <= 16'h1028	;
				14'b01111010110111: Data_out <= 16'h101B	;
				14'b01111010111000: Data_out <= 16'h100F	;
				14'b01111010111001: Data_out <= 16'h1002	;
				14'b01111010111010: Data_out <= 16'h0FF6	;
				14'b01111010111011: Data_out <= 16'h0FE9	;
				14'b01111010111100: Data_out <= 16'h0FDD	;
				14'b01111010111101: Data_out <= 16'h0FD1	;
				14'b01111010111110: Data_out <= 16'h0FC4	;
				14'b01111010111111: Data_out <= 16'h0FB8	;
				14'b01111011000000: Data_out <= 16'h0FAB	;
				14'b01111011000001: Data_out <= 16'h0F9F	;
				14'b01111011000010: Data_out <= 16'h0F92	;
				14'b01111011000011: Data_out <= 16'h0F86	;
				14'b01111011000100: Data_out <= 16'h0F79	;
				14'b01111011000101: Data_out <= 16'h0F6D	;
				14'b01111011000110: Data_out <= 16'h0F60	;
				14'b01111011000111: Data_out <= 16'h0F54	;
				14'b01111011001000: Data_out <= 16'h0F47	;
				14'b01111011001001: Data_out <= 16'h0F3B	;
				14'b01111011001010: Data_out <= 16'h0F2E	;
				14'b01111011001011: Data_out <= 16'h0F22	;
				14'b01111011001100: Data_out <= 16'h0F15	;
				14'b01111011001101: Data_out <= 16'h0F09	;
				14'b01111011001110: Data_out <= 16'h0EFC	;
				14'b01111011001111: Data_out <= 16'h0EF0	;
				14'b01111011010000: Data_out <= 16'h0EE4	;
				14'b01111011010001: Data_out <= 16'h0ED7	;
				14'b01111011010010: Data_out <= 16'h0ECB	;
				14'b01111011010011: Data_out <= 16'h0EBE	;
				14'b01111011010100: Data_out <= 16'h0EB2	;
				14'b01111011010101: Data_out <= 16'h0EA5	;
				14'b01111011010110: Data_out <= 16'h0E99	;
				14'b01111011010111: Data_out <= 16'h0E8C	;
				14'b01111011011000: Data_out <= 16'h0E80	;
				14'b01111011011001: Data_out <= 16'h0E73	;
				14'b01111011011010: Data_out <= 16'h0E67	;
				14'b01111011011011: Data_out <= 16'h0E5A	;
				14'b01111011011100: Data_out <= 16'h0E4E	;
				14'b01111011011101: Data_out <= 16'h0E41	;
				14'b01111011011110: Data_out <= 16'h0E35	;
				14'b01111011011111: Data_out <= 16'h0E28	;
				14'b01111011100000: Data_out <= 16'h0E1C	;
				14'b01111011100001: Data_out <= 16'h0E0F	;
				14'b01111011100010: Data_out <= 16'h0E03	;
				14'b01111011100011: Data_out <= 16'h0DF6	;
				14'b01111011100100: Data_out <= 16'h0DEA	;
				14'b01111011100101: Data_out <= 16'h0DDD	;
				14'b01111011100110: Data_out <= 16'h0DD1	;
				14'b01111011100111: Data_out <= 16'h0DC4	;
				14'b01111011101000: Data_out <= 16'h0DB8	;
				14'b01111011101001: Data_out <= 16'h0DAB	;
				14'b01111011101010: Data_out <= 16'h0D9F	;
				14'b01111011101011: Data_out <= 16'h0D92	;
				14'b01111011101100: Data_out <= 16'h0D86	;
				14'b01111011101101: Data_out <= 16'h0D79	;
				14'b01111011101110: Data_out <= 16'h0D6D	;
				14'b01111011101111: Data_out <= 16'h0D60	;
				14'b01111011110000: Data_out <= 16'h0D54	;
				14'b01111011110001: Data_out <= 16'h0D47	;
				14'b01111011110010: Data_out <= 16'h0D3B	;
				14'b01111011110011: Data_out <= 16'h0D2E	;
				14'b01111011110100: Data_out <= 16'h0D22	;
				14'b01111011110101: Data_out <= 16'h0D15	;
				14'b01111011110110: Data_out <= 16'h0D09	;
				14'b01111011110111: Data_out <= 16'h0CFC	;
				14'b01111011111000: Data_out <= 16'h0CF0	;
				14'b01111011111001: Data_out <= 16'h0CE3	;
				14'b01111011111010: Data_out <= 16'h0CD7	;
				14'b01111011111011: Data_out <= 16'h0CCA	;
				14'b01111011111100: Data_out <= 16'h0CBE	;
				14'b01111011111101: Data_out <= 16'h0CB1	;
				14'b01111011111110: Data_out <= 16'h0CA5	;
				14'b01111011111111: Data_out <= 16'h0C98	;
				14'b01111100000000: Data_out <= 16'h0C8C	;
				14'b01111100000001: Data_out <= 16'h0C7F	;
				14'b01111100000010: Data_out <= 16'h0C73	;
				14'b01111100000011: Data_out <= 16'h0C66	;
				14'b01111100000100: Data_out <= 16'h0C5A	;
				14'b01111100000101: Data_out <= 16'h0C4D	;
				14'b01111100000110: Data_out <= 16'h0C41	;
				14'b01111100000111: Data_out <= 16'h0C34	;
				14'b01111100001000: Data_out <= 16'h0C28	;
				14'b01111100001001: Data_out <= 16'h0C1B	;
				14'b01111100001010: Data_out <= 16'h0C0F	;
				14'b01111100001011: Data_out <= 16'h0C02	;
				14'b01111100001100: Data_out <= 16'h0BF6	;
				14'b01111100001101: Data_out <= 16'h0BE9	;
				14'b01111100001110: Data_out <= 16'h0BDD	;
				14'b01111100001111: Data_out <= 16'h0BD0	;
				14'b01111100010000: Data_out <= 16'h0BC4	;
				14'b01111100010001: Data_out <= 16'h0BB7	;
				14'b01111100010010: Data_out <= 16'h0BAB	;
				14'b01111100010011: Data_out <= 16'h0B9E	;
				14'b01111100010100: Data_out <= 16'h0B92	;
				14'b01111100010101: Data_out <= 16'h0B85	;
				14'b01111100010110: Data_out <= 16'h0B79	;
				14'b01111100010111: Data_out <= 16'h0B6C	;
				14'b01111100011000: Data_out <= 16'h0B60	;
				14'b01111100011001: Data_out <= 16'h0B53	;
				14'b01111100011010: Data_out <= 16'h0B47	;
				14'b01111100011011: Data_out <= 16'h0B3A	;
				14'b01111100011100: Data_out <= 16'h0B2D	;
				14'b01111100011101: Data_out <= 16'h0B21	;
				14'b01111100011110: Data_out <= 16'h0B14	;
				14'b01111100011111: Data_out <= 16'h0B08	;
				14'b01111100100000: Data_out <= 16'h0AFB	;
				14'b01111100100001: Data_out <= 16'h0AEF	;
				14'b01111100100010: Data_out <= 16'h0AE2	;
				14'b01111100100011: Data_out <= 16'h0AD6	;
				14'b01111100100100: Data_out <= 16'h0AC9	;
				14'b01111100100101: Data_out <= 16'h0ABD	;
				14'b01111100100110: Data_out <= 16'h0AB0	;
				14'b01111100100111: Data_out <= 16'h0AA4	;
				14'b01111100101000: Data_out <= 16'h0A97	;
				14'b01111100101001: Data_out <= 16'h0A8B	;
				14'b01111100101010: Data_out <= 16'h0A7E	;
				14'b01111100101011: Data_out <= 16'h0A72	;
				14'b01111100101100: Data_out <= 16'h0A65	;
				14'b01111100101101: Data_out <= 16'h0A59	;
				14'b01111100101110: Data_out <= 16'h0A4C	;
				14'b01111100101111: Data_out <= 16'h0A40	;
				14'b01111100110000: Data_out <= 16'h0A33	;
				14'b01111100110001: Data_out <= 16'h0A27	;
				14'b01111100110010: Data_out <= 16'h0A1A	;
				14'b01111100110011: Data_out <= 16'h0A0D	;
				14'b01111100110100: Data_out <= 16'h0A01	;
				14'b01111100110101: Data_out <= 16'h09F4	;
				14'b01111100110110: Data_out <= 16'h09E8	;
				14'b01111100110111: Data_out <= 16'h09DB	;
				14'b01111100111000: Data_out <= 16'h09CF	;
				14'b01111100111001: Data_out <= 16'h09C2	;
				14'b01111100111010: Data_out <= 16'h09B6	;
				14'b01111100111011: Data_out <= 16'h09A9	;
				14'b01111100111100: Data_out <= 16'h099D	;
				14'b01111100111101: Data_out <= 16'h0990	;
				14'b01111100111110: Data_out <= 16'h0984	;
				14'b01111100111111: Data_out <= 16'h0977	;
				14'b01111101000000: Data_out <= 16'h096B	;
				14'b01111101000001: Data_out <= 16'h095E	;
				14'b01111101000010: Data_out <= 16'h0952	;
				14'b01111101000011: Data_out <= 16'h0945	;
				14'b01111101000100: Data_out <= 16'h0938	;
				14'b01111101000101: Data_out <= 16'h092C	;
				14'b01111101000110: Data_out <= 16'h091F	;
				14'b01111101000111: Data_out <= 16'h0913	;
				14'b01111101001000: Data_out <= 16'h0906	;
				14'b01111101001001: Data_out <= 16'h08FA	;
				14'b01111101001010: Data_out <= 16'h08ED	;
				14'b01111101001011: Data_out <= 16'h08E1	;
				14'b01111101001100: Data_out <= 16'h08D4	;
				14'b01111101001101: Data_out <= 16'h08C8	;
				14'b01111101001110: Data_out <= 16'h08BB	;
				14'b01111101001111: Data_out <= 16'h08AF	;
				14'b01111101010000: Data_out <= 16'h08A2	;
				14'b01111101010001: Data_out <= 16'h0895	;
				14'b01111101010010: Data_out <= 16'h0889	;
				14'b01111101010011: Data_out <= 16'h087C	;
				14'b01111101010100: Data_out <= 16'h0870	;
				14'b01111101010101: Data_out <= 16'h0863	;
				14'b01111101010110: Data_out <= 16'h0857	;
				14'b01111101010111: Data_out <= 16'h084A	;
				14'b01111101011000: Data_out <= 16'h083E	;
				14'b01111101011001: Data_out <= 16'h0831	;
				14'b01111101011010: Data_out <= 16'h0825	;
				14'b01111101011011: Data_out <= 16'h0818	;
				14'b01111101011100: Data_out <= 16'h080C	;
				14'b01111101011101: Data_out <= 16'h07FF	;
				14'b01111101011110: Data_out <= 16'h07F2	;
				14'b01111101011111: Data_out <= 16'h07E6	;
				14'b01111101100000: Data_out <= 16'h07D9	;
				14'b01111101100001: Data_out <= 16'h07CD	;
				14'b01111101100010: Data_out <= 16'h07C0	;
				14'b01111101100011: Data_out <= 16'h07B4	;
				14'b01111101100100: Data_out <= 16'h07A7	;
				14'b01111101100101: Data_out <= 16'h079B	;
				14'b01111101100110: Data_out <= 16'h078E	;
				14'b01111101100111: Data_out <= 16'h0782	;
				14'b01111101101000: Data_out <= 16'h0775	;
				14'b01111101101001: Data_out <= 16'h0769	;
				14'b01111101101010: Data_out <= 16'h075C	;
				14'b01111101101011: Data_out <= 16'h074F	;
				14'b01111101101100: Data_out <= 16'h0743	;
				14'b01111101101101: Data_out <= 16'h0736	;
				14'b01111101101110: Data_out <= 16'h072A	;
				14'b01111101101111: Data_out <= 16'h071D	;
				14'b01111101110000: Data_out <= 16'h0711	;
				14'b01111101110001: Data_out <= 16'h0704	;
				14'b01111101110010: Data_out <= 16'h06F8	;
				14'b01111101110011: Data_out <= 16'h06EB	;
				14'b01111101110100: Data_out <= 16'h06DE	;
				14'b01111101110101: Data_out <= 16'h06D2	;
				14'b01111101110110: Data_out <= 16'h06C5	;
				14'b01111101110111: Data_out <= 16'h06B9	;
				14'b01111101111000: Data_out <= 16'h06AC	;
				14'b01111101111001: Data_out <= 16'h06A0	;
				14'b01111101111010: Data_out <= 16'h0693	;
				14'b01111101111011: Data_out <= 16'h0687	;
				14'b01111101111100: Data_out <= 16'h067A	;
				14'b01111101111101: Data_out <= 16'h066E	;
				14'b01111101111110: Data_out <= 16'h0661	;
				14'b01111101111111: Data_out <= 16'h0654	;
				14'b01111110000000: Data_out <= 16'h0648	;
				14'b01111110000001: Data_out <= 16'h063B	;
				14'b01111110000010: Data_out <= 16'h062F	;
				14'b01111110000011: Data_out <= 16'h0622	;
				14'b01111110000100: Data_out <= 16'h0616	;
				14'b01111110000101: Data_out <= 16'h0609	;
				14'b01111110000110: Data_out <= 16'h05FD	;
				14'b01111110000111: Data_out <= 16'h05F0	;
				14'b01111110001000: Data_out <= 16'h05E3	;
				14'b01111110001001: Data_out <= 16'h05D7	;
				14'b01111110001010: Data_out <= 16'h05CA	;
				14'b01111110001011: Data_out <= 16'h05BE	;
				14'b01111110001100: Data_out <= 16'h05B1	;
				14'b01111110001101: Data_out <= 16'h05A5	;
				14'b01111110001110: Data_out <= 16'h0598	;
				14'b01111110001111: Data_out <= 16'h058C	;
				14'b01111110010000: Data_out <= 16'h057F	;
				14'b01111110010001: Data_out <= 16'h0573	;
				14'b01111110010010: Data_out <= 16'h0566	;
				14'b01111110010011: Data_out <= 16'h0559	;
				14'b01111110010100: Data_out <= 16'h054D	;
				14'b01111110010101: Data_out <= 16'h0540	;
				14'b01111110010110: Data_out <= 16'h0534	;
				14'b01111110010111: Data_out <= 16'h0527	;
				14'b01111110011000: Data_out <= 16'h051B	;
				14'b01111110011001: Data_out <= 16'h050E	;
				14'b01111110011010: Data_out <= 16'h0502	;
				14'b01111110011011: Data_out <= 16'h04F5	;
				14'b01111110011100: Data_out <= 16'h04E8	;
				14'b01111110011101: Data_out <= 16'h04DC	;
				14'b01111110011110: Data_out <= 16'h04CF	;
				14'b01111110011111: Data_out <= 16'h04C3	;
				14'b01111110100000: Data_out <= 16'h04B6	;
				14'b01111110100001: Data_out <= 16'h04AA	;
				14'b01111110100010: Data_out <= 16'h049D	;
				14'b01111110100011: Data_out <= 16'h0490	;
				14'b01111110100100: Data_out <= 16'h0484	;
				14'b01111110100101: Data_out <= 16'h0477	;
				14'b01111110100110: Data_out <= 16'h046B	;
				14'b01111110100111: Data_out <= 16'h045E	;
				14'b01111110101000: Data_out <= 16'h0452	;
				14'b01111110101001: Data_out <= 16'h0445	;
				14'b01111110101010: Data_out <= 16'h0439	;
				14'b01111110101011: Data_out <= 16'h042C	;
				14'b01111110101100: Data_out <= 16'h041F	;
				14'b01111110101101: Data_out <= 16'h0413	;
				14'b01111110101110: Data_out <= 16'h0406	;
				14'b01111110101111: Data_out <= 16'h03FA	;
				14'b01111110110000: Data_out <= 16'h03ED	;
				14'b01111110110001: Data_out <= 16'h03E1	;
				14'b01111110110010: Data_out <= 16'h03D4	;
				14'b01111110110011: Data_out <= 16'h03C8	;
				14'b01111110110100: Data_out <= 16'h03BB	;
				14'b01111110110101: Data_out <= 16'h03AE	;
				14'b01111110110110: Data_out <= 16'h03A2	;
				14'b01111110110111: Data_out <= 16'h0395	;
				14'b01111110111000: Data_out <= 16'h0389	;
				14'b01111110111001: Data_out <= 16'h037C	;
				14'b01111110111010: Data_out <= 16'h0370	;
				14'b01111110111011: Data_out <= 16'h0363	;
				14'b01111110111100: Data_out <= 16'h0356	;
				14'b01111110111101: Data_out <= 16'h034A	;
				14'b01111110111110: Data_out <= 16'h033D	;
				14'b01111110111111: Data_out <= 16'h0331	;
				14'b01111111000000: Data_out <= 16'h0324	;
				14'b01111111000001: Data_out <= 16'h0318	;
				14'b01111111000010: Data_out <= 16'h030B	;
				14'b01111111000011: Data_out <= 16'h02FF	;
				14'b01111111000100: Data_out <= 16'h02F2	;
				14'b01111111000101: Data_out <= 16'h02E5	;
				14'b01111111000110: Data_out <= 16'h02D9	;
				14'b01111111000111: Data_out <= 16'h02CC	;
				14'b01111111001000: Data_out <= 16'h02C0	;
				14'b01111111001001: Data_out <= 16'h02B3	;
				14'b01111111001010: Data_out <= 16'h02A7	;
				14'b01111111001011: Data_out <= 16'h029A	;
				14'b01111111001100: Data_out <= 16'h028D	;
				14'b01111111001101: Data_out <= 16'h0281	;
				14'b01111111001110: Data_out <= 16'h0274	;
				14'b01111111001111: Data_out <= 16'h0268	;
				14'b01111111010000: Data_out <= 16'h025B	;
				14'b01111111010001: Data_out <= 16'h024F	;
				14'b01111111010010: Data_out <= 16'h0242	;
				14'b01111111010011: Data_out <= 16'h0236	;
				14'b01111111010100: Data_out <= 16'h0229	;
				14'b01111111010101: Data_out <= 16'h021C	;
				14'b01111111010110: Data_out <= 16'h0210	;
				14'b01111111010111: Data_out <= 16'h0203	;
				14'b01111111011000: Data_out <= 16'h01F7	;
				14'b01111111011001: Data_out <= 16'h01EA	;
				14'b01111111011010: Data_out <= 16'h01DE	;
				14'b01111111011011: Data_out <= 16'h01D1	;
				14'b01111111011100: Data_out <= 16'h01C4	;
				14'b01111111011101: Data_out <= 16'h01B8	;
				14'b01111111011110: Data_out <= 16'h01AB	;
				14'b01111111011111: Data_out <= 16'h019F	;
				14'b01111111100000: Data_out <= 16'h0192	;
				14'b01111111100001: Data_out <= 16'h0186	;
				14'b01111111100010: Data_out <= 16'h0179	;
				14'b01111111100011: Data_out <= 16'h016D	;
				14'b01111111100100: Data_out <= 16'h0160	;
				14'b01111111100101: Data_out <= 16'h0153	;
				14'b01111111100110: Data_out <= 16'h0147	;
				14'b01111111100111: Data_out <= 16'h013A	;
				14'b01111111101000: Data_out <= 16'h012E	;
				14'b01111111101001: Data_out <= 16'h0121	;
				14'b01111111101010: Data_out <= 16'h0115	;
				14'b01111111101011: Data_out <= 16'h0108	;
				14'b01111111101100: Data_out <= 16'h00FB	;
				14'b01111111101101: Data_out <= 16'h00EF	;
				14'b01111111101110: Data_out <= 16'h00E2	;
				14'b01111111101111: Data_out <= 16'h00D6	;
				14'b01111111110000: Data_out <= 16'h00C9	;
				14'b01111111110001: Data_out <= 16'h00BD	;
				14'b01111111110010: Data_out <= 16'h00B0	;
				14'b01111111110011: Data_out <= 16'h00A3	;
				14'b01111111110100: Data_out <= 16'h0097	;
				14'b01111111110101: Data_out <= 16'h008A	;
				14'b01111111110110: Data_out <= 16'h007E	;
				14'b01111111110111: Data_out <= 16'h0071	;
				14'b01111111111000: Data_out <= 16'h0065	;
				14'b01111111111001: Data_out <= 16'h0058	;
				14'b01111111111010: Data_out <= 16'h004B	;
				14'b01111111111011: Data_out <= 16'h003F	;
				14'b01111111111100: Data_out <= 16'h0032	;
				14'b01111111111101: Data_out <= 16'h0026	;
				14'b01111111111110: Data_out <= 16'h0019	;
				14'b01111111111111: Data_out <= 16'h000D	;
				/////////////////////////////////////////////////////////////////////////////////////////////
				//	negative	half-cycle of fall......
				14'b10000000000000: Data_out <= 16'h0000	;
				14'b10000000000001: Data_out <= 16'hFFF4	;
				14'b10000000000010: Data_out <= 16'hFFE7	;
				14'b10000000000011: Data_out <= 16'hFFDA	;
				14'b10000000000100: Data_out <= 16'hFFCE	;
				14'b10000000000101: Data_out <= 16'hFFC1	;
				14'b10000000000110: Data_out <= 16'hFFB5	;
				14'b10000000000111: Data_out <= 16'hFFA8	;
				14'b10000000001000: Data_out <= 16'hFF9C	;
				14'b10000000001001: Data_out <= 16'hFF8F	;
				14'b10000000001010: Data_out <= 16'hFF82	;
				14'b10000000001011: Data_out <= 16'hFF76	;
				14'b10000000001100: Data_out <= 16'hFF69	;
				14'b10000000001101: Data_out <= 16'hFF5D	;
				14'b10000000001110: Data_out <= 16'hFF50	;
				14'b10000000001111: Data_out <= 16'hFF44	;
				14'b10000000010000: Data_out <= 16'hFF37	;
				14'b10000000010001: Data_out <= 16'hFF2A	;
				14'b10000000010010: Data_out <= 16'hFF1E	;
				14'b10000000010011: Data_out <= 16'hFF11	;
				14'b10000000010100: Data_out <= 16'hFF05	;
				14'b10000000010101: Data_out <= 16'hFEF8	;
				14'b10000000010110: Data_out <= 16'hFEEC	;
				14'b10000000010111: Data_out <= 16'hFEDF	;
				14'b10000000011000: Data_out <= 16'hFED3	;
				14'b10000000011001: Data_out <= 16'hFEC6	;
				14'b10000000011010: Data_out <= 16'hFEB9	;
				14'b10000000011011: Data_out <= 16'hFEAD	;
				14'b10000000011100: Data_out <= 16'hFEA0	;
				14'b10000000011101: Data_out <= 16'hFE94	;
				14'b10000000011110: Data_out <= 16'hFE87	;
				14'b10000000011111: Data_out <= 16'hFE7B	;
				14'b10000000100000: Data_out <= 16'hFE6E	;
				14'b10000000100001: Data_out <= 16'hFE61	;
				14'b10000000100010: Data_out <= 16'hFE55	;
				14'b10000000100011: Data_out <= 16'hFE48	;
				14'b10000000100100: Data_out <= 16'hFE3C	;
				14'b10000000100101: Data_out <= 16'hFE2F	;
				14'b10000000100110: Data_out <= 16'hFE23	;
				14'b10000000100111: Data_out <= 16'hFE16	;
				14'b10000000101000: Data_out <= 16'hFE09	;
				14'b10000000101001: Data_out <= 16'hFDFD	;
				14'b10000000101010: Data_out <= 16'hFDF0	;
				14'b10000000101011: Data_out <= 16'hFDE4	;
				14'b10000000101100: Data_out <= 16'hFDD7	;
				14'b10000000101101: Data_out <= 16'hFDCB	;
				14'b10000000101110: Data_out <= 16'hFDBE	;
				14'b10000000101111: Data_out <= 16'hFDB2	;
				14'b10000000110000: Data_out <= 16'hFDA5	;
				14'b10000000110001: Data_out <= 16'hFD98	;
				14'b10000000110010: Data_out <= 16'hFD8C	;
				14'b10000000110011: Data_out <= 16'hFD7F	;
				14'b10000000110100: Data_out <= 16'hFD73	;
				14'b10000000110101: Data_out <= 16'hFD66	;
				14'b10000000110110: Data_out <= 16'hFD5A	;
				14'b10000000110111: Data_out <= 16'hFD4D	;
				14'b10000000111000: Data_out <= 16'hFD40	;
				14'b10000000111001: Data_out <= 16'hFD34	;
				14'b10000000111010: Data_out <= 16'hFD27	;
				14'b10000000111011: Data_out <= 16'hFD1B	;
				14'b10000000111100: Data_out <= 16'hFD0E	;
				14'b10000000111101: Data_out <= 16'hFD02	;
				14'b10000000111110: Data_out <= 16'hFCF5	;
				14'b10000000111111: Data_out <= 16'hFCE9	;
				14'b10000001000000: Data_out <= 16'hFCDC	;
				14'b10000001000001: Data_out <= 16'hFCCF	;
				14'b10000001000010: Data_out <= 16'hFCC3	;
				14'b10000001000011: Data_out <= 16'hFCB6	;
				14'b10000001000100: Data_out <= 16'hFCAA	;
				14'b10000001000101: Data_out <= 16'hFC9D	;
				14'b10000001000110: Data_out <= 16'hFC91	;
				14'b10000001000111: Data_out <= 16'hFC84	;
				14'b10000001001000: Data_out <= 16'hFC77	;
				14'b10000001001001: Data_out <= 16'hFC6B	;
				14'b10000001001010: Data_out <= 16'hFC5E	;
				14'b10000001001011: Data_out <= 16'hFC52	;
				14'b10000001001100: Data_out <= 16'hFC45	;
				14'b10000001001101: Data_out <= 16'hFC39	;
				14'b10000001001110: Data_out <= 16'hFC2C	;
				14'b10000001001111: Data_out <= 16'hFC20	;
				14'b10000001010000: Data_out <= 16'hFC13	;
				14'b10000001010001: Data_out <= 16'hFC06	;
				14'b10000001010010: Data_out <= 16'hFBFA	;
				14'b10000001010011: Data_out <= 16'hFBED	;
				14'b10000001010100: Data_out <= 16'hFBE1	;
				14'b10000001010101: Data_out <= 16'hFBD4	;
				14'b10000001010110: Data_out <= 16'hFBC8	;
				14'b10000001010111: Data_out <= 16'hFBBB	;
				14'b10000001011000: Data_out <= 16'hFBAF	;
				14'b10000001011001: Data_out <= 16'hFBA2	;
				14'b10000001011010: Data_out <= 16'hFB95	;
				14'b10000001011011: Data_out <= 16'hFB89	;
				14'b10000001011100: Data_out <= 16'hFB7C	;
				14'b10000001011101: Data_out <= 16'hFB70	;
				14'b10000001011110: Data_out <= 16'hFB63	;
				14'b10000001011111: Data_out <= 16'hFB57	;
				14'b10000001100000: Data_out <= 16'hFB4A	;
				14'b10000001100001: Data_out <= 16'hFB3D	;
				14'b10000001100010: Data_out <= 16'hFB31	;
				14'b10000001100011: Data_out <= 16'hFB24	;
				14'b10000001100100: Data_out <= 16'hFB18	;
				14'b10000001100101: Data_out <= 16'hFB0B	;
				14'b10000001100110: Data_out <= 16'hFAFF	;
				14'b10000001100111: Data_out <= 16'hFAF2	;
				14'b10000001101000: Data_out <= 16'hFAE6	;
				14'b10000001101001: Data_out <= 16'hFAD9	;
				14'b10000001101010: Data_out <= 16'hFACC	;
				14'b10000001101011: Data_out <= 16'hFAC0	;
				14'b10000001101100: Data_out <= 16'hFAB3	;
				14'b10000001101101: Data_out <= 16'hFAA7	;
				14'b10000001101110: Data_out <= 16'hFA9A	;
				14'b10000001101111: Data_out <= 16'hFA8E	;
				14'b10000001110000: Data_out <= 16'hFA81	;
				14'b10000001110001: Data_out <= 16'hFA75	;
				14'b10000001110010: Data_out <= 16'hFA68	;
				14'b10000001110011: Data_out <= 16'hFA5B	;
				14'b10000001110100: Data_out <= 16'hFA4F	;
				14'b10000001110101: Data_out <= 16'hFA42	;
				14'b10000001110110: Data_out <= 16'hFA36	;
				14'b10000001110111: Data_out <= 16'hFA29	;
				14'b10000001111000: Data_out <= 16'hFA1D	;
				14'b10000001111001: Data_out <= 16'hFA10	;
				14'b10000001111010: Data_out <= 16'hFA04	;
				14'b10000001111011: Data_out <= 16'hF9F7	;
				14'b10000001111100: Data_out <= 16'hF9EB	;
				14'b10000001111101: Data_out <= 16'hF9DE	;
				14'b10000001111110: Data_out <= 16'hF9D1	;
				14'b10000001111111: Data_out <= 16'hF9C5	;
				14'b10000010000000: Data_out <= 16'hF9B8	;
				14'b10000010000001: Data_out <= 16'hF9AC	;
				14'b10000010000010: Data_out <= 16'hF99F	;
				14'b10000010000011: Data_out <= 16'hF993	;
				14'b10000010000100: Data_out <= 16'hF986	;
				14'b10000010000101: Data_out <= 16'hF97A	;
				14'b10000010000110: Data_out <= 16'hF96D	;
				14'b10000010000111: Data_out <= 16'hF960	;
				14'b10000010001000: Data_out <= 16'hF954	;
				14'b10000010001001: Data_out <= 16'hF947	;
				14'b10000010001010: Data_out <= 16'hF93B	;
				14'b10000010001011: Data_out <= 16'hF92E	;
				14'b10000010001100: Data_out <= 16'hF922	;
				14'b10000010001101: Data_out <= 16'hF915	;
				14'b10000010001110: Data_out <= 16'hF909	;
				14'b10000010001111: Data_out <= 16'hF8FC	;
				14'b10000010010000: Data_out <= 16'hF8F0	;
				14'b10000010010001: Data_out <= 16'hF8E3	;
				14'b10000010010010: Data_out <= 16'hF8D6	;
				14'b10000010010011: Data_out <= 16'hF8CA	;
				14'b10000010010100: Data_out <= 16'hF8BD	;
				14'b10000010010101: Data_out <= 16'hF8B1	;
				14'b10000010010110: Data_out <= 16'hF8A4	;
				14'b10000010010111: Data_out <= 16'hF898	;
				14'b10000010011000: Data_out <= 16'hF88B	;
				14'b10000010011001: Data_out <= 16'hF87F	;
				14'b10000010011010: Data_out <= 16'hF872	;
				14'b10000010011011: Data_out <= 16'hF866	;
				14'b10000010011100: Data_out <= 16'hF859	;
				14'b10000010011101: Data_out <= 16'hF84C	;
				14'b10000010011110: Data_out <= 16'hF840	;
				14'b10000010011111: Data_out <= 16'hF833	;
				14'b10000010100000: Data_out <= 16'hF827	;
				14'b10000010100001: Data_out <= 16'hF81A	;
				14'b10000010100010: Data_out <= 16'hF80E	;
				14'b10000010100011: Data_out <= 16'hF801	;
				14'b10000010100100: Data_out <= 16'hF7F5	;
				14'b10000010100101: Data_out <= 16'hF7E8	;
				14'b10000010100110: Data_out <= 16'hF7DC	;
				14'b10000010100111: Data_out <= 16'hF7CF	;
				14'b10000010101000: Data_out <= 16'hF7C2	;
				14'b10000010101001: Data_out <= 16'hF7B6	;
				14'b10000010101010: Data_out <= 16'hF7A9	;
				14'b10000010101011: Data_out <= 16'hF79D	;
				14'b10000010101100: Data_out <= 16'hF790	;
				14'b10000010101101: Data_out <= 16'hF784	;
				14'b10000010101110: Data_out <= 16'hF777	;
				14'b10000010101111: Data_out <= 16'hF76B	;
				14'b10000010110000: Data_out <= 16'hF75E	;
				14'b10000010110001: Data_out <= 16'hF752	;
				14'b10000010110010: Data_out <= 16'hF745	;
				14'b10000010110011: Data_out <= 16'hF739	;
				14'b10000010110100: Data_out <= 16'hF72C	;
				14'b10000010110101: Data_out <= 16'hF71F	;
				14'b10000010110110: Data_out <= 16'hF713	;
				14'b10000010110111: Data_out <= 16'hF706	;
				14'b10000010111000: Data_out <= 16'hF6FA	;
				14'b10000010111001: Data_out <= 16'hF6ED	;
				14'b10000010111010: Data_out <= 16'hF6E1	;
				14'b10000010111011: Data_out <= 16'hF6D4	;
				14'b10000010111100: Data_out <= 16'hF6C8	;
				14'b10000010111101: Data_out <= 16'hF6BB	;
				14'b10000010111110: Data_out <= 16'hF6AF	;
				14'b10000010111111: Data_out <= 16'hF6A2	;
				14'b10000011000000: Data_out <= 16'hF696	;
				14'b10000011000001: Data_out <= 16'hF689	;
				14'b10000011000010: Data_out <= 16'hF67D	;
				14'b10000011000011: Data_out <= 16'hF670	;
				14'b10000011000100: Data_out <= 16'hF663	;
				14'b10000011000101: Data_out <= 16'hF657	;
				14'b10000011000110: Data_out <= 16'hF64A	;
				14'b10000011000111: Data_out <= 16'hF63E	;
				14'b10000011001000: Data_out <= 16'hF631	;
				14'b10000011001001: Data_out <= 16'hF625	;
				14'b10000011001010: Data_out <= 16'hF618	;
				14'b10000011001011: Data_out <= 16'hF60C	;
				14'b10000011001100: Data_out <= 16'hF5FF	;
				14'b10000011001101: Data_out <= 16'hF5F3	;
				14'b10000011001110: Data_out <= 16'hF5E6	;
				14'b10000011001111: Data_out <= 16'hF5DA	;
				14'b10000011010000: Data_out <= 16'hF5CD	;
				14'b10000011010001: Data_out <= 16'hF5C1	;
				14'b10000011010010: Data_out <= 16'hF5B4	;
				14'b10000011010011: Data_out <= 16'hF5A8	;
				14'b10000011010100: Data_out <= 16'hF59B	;
				14'b10000011010101: Data_out <= 16'hF58F	;
				14'b10000011010110: Data_out <= 16'hF582	;
				14'b10000011010111: Data_out <= 16'hF575	;
				14'b10000011011000: Data_out <= 16'hF569	;
				14'b10000011011001: Data_out <= 16'hF55C	;
				14'b10000011011010: Data_out <= 16'hF550	;
				14'b10000011011011: Data_out <= 16'hF543	;
				14'b10000011011100: Data_out <= 16'hF537	;
				14'b10000011011101: Data_out <= 16'hF52A	;
				14'b10000011011110: Data_out <= 16'hF51E	;
				14'b10000011011111: Data_out <= 16'hF511	;
				14'b10000011100000: Data_out <= 16'hF505	;
				14'b10000011100001: Data_out <= 16'hF4F8	;
				14'b10000011100010: Data_out <= 16'hF4EC	;
				14'b10000011100011: Data_out <= 16'hF4DF	;
				14'b10000011100100: Data_out <= 16'hF4D3	;
				14'b10000011100101: Data_out <= 16'hF4C6	;
				14'b10000011100110: Data_out <= 16'hF4BA	;
				14'b10000011100111: Data_out <= 16'hF4AD	;
				14'b10000011101000: Data_out <= 16'hF4A1	;
				14'b10000011101001: Data_out <= 16'hF494	;
				14'b10000011101010: Data_out <= 16'hF488	;
				14'b10000011101011: Data_out <= 16'hF47B	;
				14'b10000011101100: Data_out <= 16'hF46F	;
				14'b10000011101101: Data_out <= 16'hF462	;
				14'b10000011101110: Data_out <= 16'hF456	;
				14'b10000011101111: Data_out <= 16'hF449	;
				14'b10000011110000: Data_out <= 16'hF43D	;
				14'b10000011110001: Data_out <= 16'hF430	;
				14'b10000011110010: Data_out <= 16'hF423	;
				14'b10000011110011: Data_out <= 16'hF417	;
				14'b10000011110100: Data_out <= 16'hF40A	;
				14'b10000011110101: Data_out <= 16'hF3FE	;
				14'b10000011110110: Data_out <= 16'hF3F1	;
				14'b10000011110111: Data_out <= 16'hF3E5	;
				14'b10000011111000: Data_out <= 16'hF3D8	;
				14'b10000011111001: Data_out <= 16'hF3CC	;
				14'b10000011111010: Data_out <= 16'hF3BF	;
				14'b10000011111011: Data_out <= 16'hF3B3	;
				14'b10000011111100: Data_out <= 16'hF3A6	;
				14'b10000011111101: Data_out <= 16'hF39A	;
				14'b10000011111110: Data_out <= 16'hF38D	;
				14'b10000011111111: Data_out <= 16'hF381	;
				14'b10000100000000: Data_out <= 16'hF374	;
				14'b10000100000001: Data_out <= 16'hF368	;
				14'b10000100000010: Data_out <= 16'hF35B	;
				14'b10000100000011: Data_out <= 16'hF34F	;
				14'b10000100000100: Data_out <= 16'hF342	;
				14'b10000100000101: Data_out <= 16'hF336	;
				14'b10000100000110: Data_out <= 16'hF329	;
				14'b10000100000111: Data_out <= 16'hF31D	;
				14'b10000100001000: Data_out <= 16'hF310	;
				14'b10000100001001: Data_out <= 16'hF304	;
				14'b10000100001010: Data_out <= 16'hF2F7	;
				14'b10000100001011: Data_out <= 16'hF2EB	;
				14'b10000100001100: Data_out <= 16'hF2DE	;
				14'b10000100001101: Data_out <= 16'hF2D2	;
				14'b10000100001110: Data_out <= 16'hF2C5	;
				14'b10000100001111: Data_out <= 16'hF2B9	;
				14'b10000100010000: Data_out <= 16'hF2AC	;
				14'b10000100010001: Data_out <= 16'hF2A0	;
				14'b10000100010010: Data_out <= 16'hF293	;
				14'b10000100010011: Data_out <= 16'hF287	;
				14'b10000100010100: Data_out <= 16'hF27A	;
				14'b10000100010101: Data_out <= 16'hF26E	;
				14'b10000100010110: Data_out <= 16'hF261	;
				14'b10000100010111: Data_out <= 16'hF255	;
				14'b10000100011000: Data_out <= 16'hF248	;
				14'b10000100011001: Data_out <= 16'hF23C	;
				14'b10000100011010: Data_out <= 16'hF22F	;
				14'b10000100011011: Data_out <= 16'hF223	;
				14'b10000100011100: Data_out <= 16'hF216	;
				14'b10000100011101: Data_out <= 16'hF20A	;
				14'b10000100011110: Data_out <= 16'hF1FD	;
				14'b10000100011111: Data_out <= 16'hF1F1	;
				14'b10000100100000: Data_out <= 16'hF1E4	;
				14'b10000100100001: Data_out <= 16'hF1D8	;
				14'b10000100100010: Data_out <= 16'hF1CB	;
				14'b10000100100011: Data_out <= 16'hF1BF	;
				14'b10000100100100: Data_out <= 16'hF1B2	;
				14'b10000100100101: Data_out <= 16'hF1A6	;
				14'b10000100100110: Data_out <= 16'hF19A	;
				14'b10000100100111: Data_out <= 16'hF18D	;
				14'b10000100101000: Data_out <= 16'hF181	;
				14'b10000100101001: Data_out <= 16'hF174	;
				14'b10000100101010: Data_out <= 16'hF168	;
				14'b10000100101011: Data_out <= 16'hF15B	;
				14'b10000100101100: Data_out <= 16'hF14F	;
				14'b10000100101101: Data_out <= 16'hF142	;
				14'b10000100101110: Data_out <= 16'hF136	;
				14'b10000100101111: Data_out <= 16'hF129	;
				14'b10000100110000: Data_out <= 16'hF11D	;
				14'b10000100110001: Data_out <= 16'hF110	;
				14'b10000100110010: Data_out <= 16'hF104	;
				14'b10000100110011: Data_out <= 16'hF0F7	;
				14'b10000100110100: Data_out <= 16'hF0EB	;
				14'b10000100110101: Data_out <= 16'hF0DE	;
				14'b10000100110110: Data_out <= 16'hF0D2	;
				14'b10000100110111: Data_out <= 16'hF0C5	;
				14'b10000100111000: Data_out <= 16'hF0B9	;
				14'b10000100111001: Data_out <= 16'hF0AC	;
				14'b10000100111010: Data_out <= 16'hF0A0	;
				14'b10000100111011: Data_out <= 16'hF093	;
				14'b10000100111100: Data_out <= 16'hF087	;
				14'b10000100111101: Data_out <= 16'hF07A	;
				14'b10000100111110: Data_out <= 16'hF06E	;
				14'b10000100111111: Data_out <= 16'hF062	;
				14'b10000101000000: Data_out <= 16'hF055	;
				14'b10000101000001: Data_out <= 16'hF049	;
				14'b10000101000010: Data_out <= 16'hF03C	;
				14'b10000101000011: Data_out <= 16'hF030	;
				14'b10000101000100: Data_out <= 16'hF023	;
				14'b10000101000101: Data_out <= 16'hF017	;
				14'b10000101000110: Data_out <= 16'hF00A	;
				14'b10000101000111: Data_out <= 16'hEFFE	;
				14'b10000101001000: Data_out <= 16'hEFF1	;
				14'b10000101001001: Data_out <= 16'hEFE5	;
				14'b10000101001010: Data_out <= 16'hEFD8	;
				14'b10000101001011: Data_out <= 16'hEFCC	;
				14'b10000101001100: Data_out <= 16'hEFBF	;
				14'b10000101001101: Data_out <= 16'hEFB3	;
				14'b10000101001110: Data_out <= 16'hEFA7	;
				14'b10000101001111: Data_out <= 16'hEF9A	;
				14'b10000101010000: Data_out <= 16'hEF8E	;
				14'b10000101010001: Data_out <= 16'hEF81	;
				14'b10000101010010: Data_out <= 16'hEF75	;
				14'b10000101010011: Data_out <= 16'hEF68	;
				14'b10000101010100: Data_out <= 16'hEF5C	;
				14'b10000101010101: Data_out <= 16'hEF4F	;
				14'b10000101010110: Data_out <= 16'hEF43	;
				14'b10000101010111: Data_out <= 16'hEF36	;
				14'b10000101011000: Data_out <= 16'hEF2A	;
				14'b10000101011001: Data_out <= 16'hEF1D	;
				14'b10000101011010: Data_out <= 16'hEF11	;
				14'b10000101011011: Data_out <= 16'hEF05	;
				14'b10000101011100: Data_out <= 16'hEEF8	;
				14'b10000101011101: Data_out <= 16'hEEEC	;
				14'b10000101011110: Data_out <= 16'hEEDF	;
				14'b10000101011111: Data_out <= 16'hEED3	;
				14'b10000101100000: Data_out <= 16'hEEC6	;
				14'b10000101100001: Data_out <= 16'hEEBA	;
				14'b10000101100010: Data_out <= 16'hEEAD	;
				14'b10000101100011: Data_out <= 16'hEEA1	;
				14'b10000101100100: Data_out <= 16'hEE94	;
				14'b10000101100101: Data_out <= 16'hEE88	;
				14'b10000101100110: Data_out <= 16'hEE7C	;
				14'b10000101100111: Data_out <= 16'hEE6F	;
				14'b10000101101000: Data_out <= 16'hEE63	;
				14'b10000101101001: Data_out <= 16'hEE56	;
				14'b10000101101010: Data_out <= 16'hEE4A	;
				14'b10000101101011: Data_out <= 16'hEE3D	;
				14'b10000101101100: Data_out <= 16'hEE31	;
				14'b10000101101101: Data_out <= 16'hEE24	;
				14'b10000101101110: Data_out <= 16'hEE18	;
				14'b10000101101111: Data_out <= 16'hEE0C	;
				14'b10000101110000: Data_out <= 16'hEDFF	;
				14'b10000101110001: Data_out <= 16'hEDF3	;
				14'b10000101110010: Data_out <= 16'hEDE6	;
				14'b10000101110011: Data_out <= 16'hEDDA	;
				14'b10000101110100: Data_out <= 16'hEDCD	;
				14'b10000101110101: Data_out <= 16'hEDC1	;
				14'b10000101110110: Data_out <= 16'hEDB5	;
				14'b10000101110111: Data_out <= 16'hEDA8	;
				14'b10000101111000: Data_out <= 16'hED9C	;
				14'b10000101111001: Data_out <= 16'hED8F	;
				14'b10000101111010: Data_out <= 16'hED83	;
				14'b10000101111011: Data_out <= 16'hED76	;
				14'b10000101111100: Data_out <= 16'hED6A	;
				14'b10000101111101: Data_out <= 16'hED5D	;
				14'b10000101111110: Data_out <= 16'hED51	;
				14'b10000101111111: Data_out <= 16'hED45	;
				14'b10000110000000: Data_out <= 16'hED38	;
				14'b10000110000001: Data_out <= 16'hED2C	;
				14'b10000110000010: Data_out <= 16'hED1F	;
				14'b10000110000011: Data_out <= 16'hED13	;
				14'b10000110000100: Data_out <= 16'hED06	;
				14'b10000110000101: Data_out <= 16'hECFA	;
				14'b10000110000110: Data_out <= 16'hECEE	;
				14'b10000110000111: Data_out <= 16'hECE1	;
				14'b10000110001000: Data_out <= 16'hECD5	;
				14'b10000110001001: Data_out <= 16'hECC8	;
				14'b10000110001010: Data_out <= 16'hECBC	;
				14'b10000110001011: Data_out <= 16'hECAF	;
				14'b10000110001100: Data_out <= 16'hECA3	;
				14'b10000110001101: Data_out <= 16'hEC97	;
				14'b10000110001110: Data_out <= 16'hEC8A	;
				14'b10000110001111: Data_out <= 16'hEC7E	;
				14'b10000110010000: Data_out <= 16'hEC71	;
				14'b10000110010001: Data_out <= 16'hEC65	;
				14'b10000110010010: Data_out <= 16'hEC59	;
				14'b10000110010011: Data_out <= 16'hEC4C	;
				14'b10000110010100: Data_out <= 16'hEC40	;
				14'b10000110010101: Data_out <= 16'hEC33	;
				14'b10000110010110: Data_out <= 16'hEC27	;
				14'b10000110010111: Data_out <= 16'hEC1A	;
				14'b10000110011000: Data_out <= 16'hEC0E	;
				14'b10000110011001: Data_out <= 16'hEC02	;
				14'b10000110011010: Data_out <= 16'hEBF5	;
				14'b10000110011011: Data_out <= 16'hEBE9	;
				14'b10000110011100: Data_out <= 16'hEBDC	;
				14'b10000110011101: Data_out <= 16'hEBD0	;
				14'b10000110011110: Data_out <= 16'hEBC4	;
				14'b10000110011111: Data_out <= 16'hEBB7	;
				14'b10000110100000: Data_out <= 16'hEBAB	;
				14'b10000110100001: Data_out <= 16'hEB9E	;
				14'b10000110100010: Data_out <= 16'hEB92	;
				14'b10000110100011: Data_out <= 16'hEB86	;
				14'b10000110100100: Data_out <= 16'hEB79	;
				14'b10000110100101: Data_out <= 16'hEB6D	;
				14'b10000110100110: Data_out <= 16'hEB60	;
				14'b10000110100111: Data_out <= 16'hEB54	;
				14'b10000110101000: Data_out <= 16'hEB48	;
				14'b10000110101001: Data_out <= 16'hEB3B	;
				14'b10000110101010: Data_out <= 16'hEB2F	;
				14'b10000110101011: Data_out <= 16'hEB22	;
				14'b10000110101100: Data_out <= 16'hEB16	;
				14'b10000110101101: Data_out <= 16'hEB0A	;
				14'b10000110101110: Data_out <= 16'hEAFD	;
				14'b10000110101111: Data_out <= 16'hEAF1	;
				14'b10000110110000: Data_out <= 16'hEAE4	;
				14'b10000110110001: Data_out <= 16'hEAD8	;
				14'b10000110110010: Data_out <= 16'hEACC	;
				14'b10000110110011: Data_out <= 16'hEABF	;
				14'b10000110110100: Data_out <= 16'hEAB3	;
				14'b10000110110101: Data_out <= 16'hEAA6	;
				14'b10000110110110: Data_out <= 16'hEA9A	;
				14'b10000110110111: Data_out <= 16'hEA8E	;
				14'b10000110111000: Data_out <= 16'hEA81	;
				14'b10000110111001: Data_out <= 16'hEA75	;
				14'b10000110111010: Data_out <= 16'hEA68	;
				14'b10000110111011: Data_out <= 16'hEA5C	;
				14'b10000110111100: Data_out <= 16'hEA50	;
				14'b10000110111101: Data_out <= 16'hEA43	;
				14'b10000110111110: Data_out <= 16'hEA37	;
				14'b10000110111111: Data_out <= 16'hEA2B	;
				14'b10000111000000: Data_out <= 16'hEA1E	;
				14'b10000111000001: Data_out <= 16'hEA12	;
				14'b10000111000010: Data_out <= 16'hEA05	;
				14'b10000111000011: Data_out <= 16'hE9F9	;
				14'b10000111000100: Data_out <= 16'hE9ED	;
				14'b10000111000101: Data_out <= 16'hE9E0	;
				14'b10000111000110: Data_out <= 16'hE9D4	;
				14'b10000111000111: Data_out <= 16'hE9C8	;
				14'b10000111001000: Data_out <= 16'hE9BB	;
				14'b10000111001001: Data_out <= 16'hE9AF	;
				14'b10000111001010: Data_out <= 16'hE9A2	;
				14'b10000111001011: Data_out <= 16'hE996	;
				14'b10000111001100: Data_out <= 16'hE98A	;
				14'b10000111001101: Data_out <= 16'hE97D	;
				14'b10000111001110: Data_out <= 16'hE971	;
				14'b10000111001111: Data_out <= 16'hE965	;
				14'b10000111010000: Data_out <= 16'hE958	;
				14'b10000111010001: Data_out <= 16'hE94C	;
				14'b10000111010010: Data_out <= 16'hE93F	;
				14'b10000111010011: Data_out <= 16'hE933	;
				14'b10000111010100: Data_out <= 16'hE927	;
				14'b10000111010101: Data_out <= 16'hE91A	;
				14'b10000111010110: Data_out <= 16'hE90E	;
				14'b10000111010111: Data_out <= 16'hE902	;
				14'b10000111011000: Data_out <= 16'hE8F5	;
				14'b10000111011001: Data_out <= 16'hE8E9	;
				14'b10000111011010: Data_out <= 16'hE8DD	;
				14'b10000111011011: Data_out <= 16'hE8D0	;
				14'b10000111011100: Data_out <= 16'hE8C4	;
				14'b10000111011101: Data_out <= 16'hE8B7	;
				14'b10000111011110: Data_out <= 16'hE8AB	;
				14'b10000111011111: Data_out <= 16'hE89F	;
				14'b10000111100000: Data_out <= 16'hE892	;
				14'b10000111100001: Data_out <= 16'hE886	;
				14'b10000111100010: Data_out <= 16'hE87A	;
				14'b10000111100011: Data_out <= 16'hE86D	;
				14'b10000111100100: Data_out <= 16'hE861	;
				14'b10000111100101: Data_out <= 16'hE855	;
				14'b10000111100110: Data_out <= 16'hE848	;
				14'b10000111100111: Data_out <= 16'hE83C	;
				14'b10000111101000: Data_out <= 16'hE830	;
				14'b10000111101001: Data_out <= 16'hE823	;
				14'b10000111101010: Data_out <= 16'hE817	;
				14'b10000111101011: Data_out <= 16'hE80B	;
				14'b10000111101100: Data_out <= 16'hE7FE	;
				14'b10000111101101: Data_out <= 16'hE7F2	;
				14'b10000111101110: Data_out <= 16'hE7E6	;
				14'b10000111101111: Data_out <= 16'hE7D9	;
				14'b10000111110000: Data_out <= 16'hE7CD	;
				14'b10000111110001: Data_out <= 16'hE7C1	;
				14'b10000111110010: Data_out <= 16'hE7B4	;
				14'b10000111110011: Data_out <= 16'hE7A8	;
				14'b10000111110100: Data_out <= 16'hE79C	;
				14'b10000111110101: Data_out <= 16'hE78F	;
				14'b10000111110110: Data_out <= 16'hE783	;
				14'b10000111110111: Data_out <= 16'hE777	;
				14'b10000111111000: Data_out <= 16'hE76A	;
				14'b10000111111001: Data_out <= 16'hE75E	;
				14'b10000111111010: Data_out <= 16'hE752	;
				14'b10000111111011: Data_out <= 16'hE745	;
				14'b10000111111100: Data_out <= 16'hE739	;
				14'b10000111111101: Data_out <= 16'hE72D	;
				14'b10000111111110: Data_out <= 16'hE720	;
				14'b10000111111111: Data_out <= 16'hE714	;
				14'b10001000000000: Data_out <= 16'hE708	;
				14'b10001000000001: Data_out <= 16'hE6FB	;
				14'b10001000000010: Data_out <= 16'hE6EF	;
				14'b10001000000011: Data_out <= 16'hE6E3	;
				14'b10001000000100: Data_out <= 16'hE6D6	;
				14'b10001000000101: Data_out <= 16'hE6CA	;
				14'b10001000000110: Data_out <= 16'hE6BE	;
				14'b10001000000111: Data_out <= 16'hE6B1	;
				14'b10001000001000: Data_out <= 16'hE6A5	;
				14'b10001000001001: Data_out <= 16'hE699	;
				14'b10001000001010: Data_out <= 16'hE68C	;
				14'b10001000001011: Data_out <= 16'hE680	;
				14'b10001000001100: Data_out <= 16'hE674	;
				14'b10001000001101: Data_out <= 16'hE667	;
				14'b10001000001110: Data_out <= 16'hE65B	;
				14'b10001000001111: Data_out <= 16'hE64F	;
				14'b10001000010000: Data_out <= 16'hE643	;
				14'b10001000010001: Data_out <= 16'hE636	;
				14'b10001000010010: Data_out <= 16'hE62A	;
				14'b10001000010011: Data_out <= 16'hE61E	;
				14'b10001000010100: Data_out <= 16'hE611	;
				14'b10001000010101: Data_out <= 16'hE605	;
				14'b10001000010110: Data_out <= 16'hE5F9	;
				14'b10001000010111: Data_out <= 16'hE5EC	;
				14'b10001000011000: Data_out <= 16'hE5E0	;
				14'b10001000011001: Data_out <= 16'hE5D4	;
				14'b10001000011010: Data_out <= 16'hE5C7	;
				14'b10001000011011: Data_out <= 16'hE5BB	;
				14'b10001000011100: Data_out <= 16'hE5AF	;
				14'b10001000011101: Data_out <= 16'hE5A3	;
				14'b10001000011110: Data_out <= 16'hE596	;
				14'b10001000011111: Data_out <= 16'hE58A	;
				14'b10001000100000: Data_out <= 16'hE57E	;
				14'b10001000100001: Data_out <= 16'hE571	;
				14'b10001000100010: Data_out <= 16'hE565	;
				14'b10001000100011: Data_out <= 16'hE559	;
				14'b10001000100100: Data_out <= 16'hE54D	;
				14'b10001000100101: Data_out <= 16'hE540	;
				14'b10001000100110: Data_out <= 16'hE534	;
				14'b10001000100111: Data_out <= 16'hE528	;
				14'b10001000101000: Data_out <= 16'hE51B	;
				14'b10001000101001: Data_out <= 16'hE50F	;
				14'b10001000101010: Data_out <= 16'hE503	;
				14'b10001000101011: Data_out <= 16'hE4F7	;
				14'b10001000101100: Data_out <= 16'hE4EA	;
				14'b10001000101101: Data_out <= 16'hE4DE	;
				14'b10001000101110: Data_out <= 16'hE4D2	;
				14'b10001000101111: Data_out <= 16'hE4C5	;
				14'b10001000110000: Data_out <= 16'hE4B9	;
				14'b10001000110001: Data_out <= 16'hE4AD	;
				14'b10001000110010: Data_out <= 16'hE4A1	;
				14'b10001000110011: Data_out <= 16'hE494	;
				14'b10001000110100: Data_out <= 16'hE488	;
				14'b10001000110101: Data_out <= 16'hE47C	;
				14'b10001000110110: Data_out <= 16'hE46F	;
				14'b10001000110111: Data_out <= 16'hE463	;
				14'b10001000111000: Data_out <= 16'hE457	;
				14'b10001000111001: Data_out <= 16'hE44B	;
				14'b10001000111010: Data_out <= 16'hE43E	;
				14'b10001000111011: Data_out <= 16'hE432	;
				14'b10001000111100: Data_out <= 16'hE426	;
				14'b10001000111101: Data_out <= 16'hE41A	;
				14'b10001000111110: Data_out <= 16'hE40D	;
				14'b10001000111111: Data_out <= 16'hE401	;
				14'b10001001000000: Data_out <= 16'hE3F5	;
				14'b10001001000001: Data_out <= 16'hE3E9	;
				14'b10001001000010: Data_out <= 16'hE3DC	;
				14'b10001001000011: Data_out <= 16'hE3D0	;
				14'b10001001000100: Data_out <= 16'hE3C4	;
				14'b10001001000101: Data_out <= 16'hE3B8	;
				14'b10001001000110: Data_out <= 16'hE3AB	;
				14'b10001001000111: Data_out <= 16'hE39F	;
				14'b10001001001000: Data_out <= 16'hE393	;
				14'b10001001001001: Data_out <= 16'hE387	;
				14'b10001001001010: Data_out <= 16'hE37A	;
				14'b10001001001011: Data_out <= 16'hE36E	;
				14'b10001001001100: Data_out <= 16'hE362	;
				14'b10001001001101: Data_out <= 16'hE356	;
				14'b10001001001110: Data_out <= 16'hE349	;
				14'b10001001001111: Data_out <= 16'hE33D	;
				14'b10001001010000: Data_out <= 16'hE331	;
				14'b10001001010001: Data_out <= 16'hE325	;
				14'b10001001010010: Data_out <= 16'hE318	;
				14'b10001001010011: Data_out <= 16'hE30C	;
				14'b10001001010100: Data_out <= 16'hE300	;
				14'b10001001010101: Data_out <= 16'hE2F4	;
				14'b10001001010110: Data_out <= 16'hE2E7	;
				14'b10001001010111: Data_out <= 16'hE2DB	;
				14'b10001001011000: Data_out <= 16'hE2CF	;
				14'b10001001011001: Data_out <= 16'hE2C3	;
				14'b10001001011010: Data_out <= 16'hE2B6	;
				14'b10001001011011: Data_out <= 16'hE2AA	;
				14'b10001001011100: Data_out <= 16'hE29E	;
				14'b10001001011101: Data_out <= 16'hE292	;
				14'b10001001011110: Data_out <= 16'hE285	;
				14'b10001001011111: Data_out <= 16'hE279	;
				14'b10001001100000: Data_out <= 16'hE26D	;
				14'b10001001100001: Data_out <= 16'hE261	;
				14'b10001001100010: Data_out <= 16'hE255	;
				14'b10001001100011: Data_out <= 16'hE248	;
				14'b10001001100100: Data_out <= 16'hE23C	;
				14'b10001001100101: Data_out <= 16'hE230	;
				14'b10001001100110: Data_out <= 16'hE224	;
				14'b10001001100111: Data_out <= 16'hE217	;
				14'b10001001101000: Data_out <= 16'hE20B	;
				14'b10001001101001: Data_out <= 16'hE1FF	;
				14'b10001001101010: Data_out <= 16'hE1F3	;
				14'b10001001101011: Data_out <= 16'hE1E7	;
				14'b10001001101100: Data_out <= 16'hE1DA	;
				14'b10001001101101: Data_out <= 16'hE1CE	;
				14'b10001001101110: Data_out <= 16'hE1C2	;
				14'b10001001101111: Data_out <= 16'hE1B6	;
				14'b10001001110000: Data_out <= 16'hE1AA	;
				14'b10001001110001: Data_out <= 16'hE19D	;
				14'b10001001110010: Data_out <= 16'hE191	;
				14'b10001001110011: Data_out <= 16'hE185	;
				14'b10001001110100: Data_out <= 16'hE179	;
				14'b10001001110101: Data_out <= 16'hE16D	;
				14'b10001001110110: Data_out <= 16'hE160	;
				14'b10001001110111: Data_out <= 16'hE154	;
				14'b10001001111000: Data_out <= 16'hE148	;
				14'b10001001111001: Data_out <= 16'hE13C	;
				14'b10001001111010: Data_out <= 16'hE130	;
				14'b10001001111011: Data_out <= 16'hE123	;
				14'b10001001111100: Data_out <= 16'hE117	;
				14'b10001001111101: Data_out <= 16'hE10B	;
				14'b10001001111110: Data_out <= 16'hE0FF	;
				14'b10001001111111: Data_out <= 16'hE0F3	;
				14'b10001010000000: Data_out <= 16'hE0E6	;
				14'b10001010000001: Data_out <= 16'hE0DA	;
				14'b10001010000010: Data_out <= 16'hE0CE	;
				14'b10001010000011: Data_out <= 16'hE0C2	;
				14'b10001010000100: Data_out <= 16'hE0B6	;
				14'b10001010000101: Data_out <= 16'hE0A9	;
				14'b10001010000110: Data_out <= 16'hE09D	;
				14'b10001010000111: Data_out <= 16'hE091	;
				14'b10001010001000: Data_out <= 16'hE085	;
				14'b10001010001001: Data_out <= 16'hE079	;
				14'b10001010001010: Data_out <= 16'hE06D	;
				14'b10001010001011: Data_out <= 16'hE060	;
				14'b10001010001100: Data_out <= 16'hE054	;
				14'b10001010001101: Data_out <= 16'hE048	;
				14'b10001010001110: Data_out <= 16'hE03C	;
				14'b10001010001111: Data_out <= 16'hE030	;
				14'b10001010010000: Data_out <= 16'hE023	;
				14'b10001010010001: Data_out <= 16'hE017	;
				14'b10001010010010: Data_out <= 16'hE00B	;
				14'b10001010010011: Data_out <= 16'hDFFF	;
				14'b10001010010100: Data_out <= 16'hDFF3	;
				14'b10001010010101: Data_out <= 16'hDFE7	;
				14'b10001010010110: Data_out <= 16'hDFDA	;
				14'b10001010010111: Data_out <= 16'hDFCE	;
				14'b10001010011000: Data_out <= 16'hDFC2	;
				14'b10001010011001: Data_out <= 16'hDFB6	;
				14'b10001010011010: Data_out <= 16'hDFAA	;
				14'b10001010011011: Data_out <= 16'hDF9E	;
				14'b10001010011100: Data_out <= 16'hDF92	;
				14'b10001010011101: Data_out <= 16'hDF85	;
				14'b10001010011110: Data_out <= 16'hDF79	;
				14'b10001010011111: Data_out <= 16'hDF6D	;
				14'b10001010100000: Data_out <= 16'hDF61	;
				14'b10001010100001: Data_out <= 16'hDF55	;
				14'b10001010100010: Data_out <= 16'hDF49	;
				14'b10001010100011: Data_out <= 16'hDF3C	;
				14'b10001010100100: Data_out <= 16'hDF30	;
				14'b10001010100101: Data_out <= 16'hDF24	;
				14'b10001010100110: Data_out <= 16'hDF18	;
				14'b10001010100111: Data_out <= 16'hDF0C	;
				14'b10001010101000: Data_out <= 16'hDF00	;
				14'b10001010101001: Data_out <= 16'hDEF4	;
				14'b10001010101010: Data_out <= 16'hDEE7	;
				14'b10001010101011: Data_out <= 16'hDEDB	;
				14'b10001010101100: Data_out <= 16'hDECF	;
				14'b10001010101101: Data_out <= 16'hDEC3	;
				14'b10001010101110: Data_out <= 16'hDEB7	;
				14'b10001010101111: Data_out <= 16'hDEAB	;
				14'b10001010110000: Data_out <= 16'hDE9F	;
				14'b10001010110001: Data_out <= 16'hDE93	;
				14'b10001010110010: Data_out <= 16'hDE86	;
				14'b10001010110011: Data_out <= 16'hDE7A	;
				14'b10001010110100: Data_out <= 16'hDE6E	;
				14'b10001010110101: Data_out <= 16'hDE62	;
				14'b10001010110110: Data_out <= 16'hDE56	;
				14'b10001010110111: Data_out <= 16'hDE4A	;
				14'b10001010111000: Data_out <= 16'hDE3E	;
				14'b10001010111001: Data_out <= 16'hDE32	;
				14'b10001010111010: Data_out <= 16'hDE25	;
				14'b10001010111011: Data_out <= 16'hDE19	;
				14'b10001010111100: Data_out <= 16'hDE0D	;
				14'b10001010111101: Data_out <= 16'hDE01	;
				14'b10001010111110: Data_out <= 16'hDDF5	;
				14'b10001010111111: Data_out <= 16'hDDE9	;
				14'b10001011000000: Data_out <= 16'hDDDD	;
				14'b10001011000001: Data_out <= 16'hDDD1	;
				14'b10001011000010: Data_out <= 16'hDDC5	;
				14'b10001011000011: Data_out <= 16'hDDB8	;
				14'b10001011000100: Data_out <= 16'hDDAC	;
				14'b10001011000101: Data_out <= 16'hDDA0	;
				14'b10001011000110: Data_out <= 16'hDD94	;
				14'b10001011000111: Data_out <= 16'hDD88	;
				14'b10001011001000: Data_out <= 16'hDD7C	;
				14'b10001011001001: Data_out <= 16'hDD70	;
				14'b10001011001010: Data_out <= 16'hDD64	;
				14'b10001011001011: Data_out <= 16'hDD58	;
				14'b10001011001100: Data_out <= 16'hDD4B	;
				14'b10001011001101: Data_out <= 16'hDD3F	;
				14'b10001011001110: Data_out <= 16'hDD33	;
				14'b10001011001111: Data_out <= 16'hDD27	;
				14'b10001011010000: Data_out <= 16'hDD1B	;
				14'b10001011010001: Data_out <= 16'hDD0F	;
				14'b10001011010010: Data_out <= 16'hDD03	;
				14'b10001011010011: Data_out <= 16'hDCF7	;
				14'b10001011010100: Data_out <= 16'hDCEB	;
				14'b10001011010101: Data_out <= 16'hDCDF	;
				14'b10001011010110: Data_out <= 16'hDCD3	;
				14'b10001011010111: Data_out <= 16'hDCC7	;
				14'b10001011011000: Data_out <= 16'hDCBA	;
				14'b10001011011001: Data_out <= 16'hDCAE	;
				14'b10001011011010: Data_out <= 16'hDCA2	;
				14'b10001011011011: Data_out <= 16'hDC96	;
				14'b10001011011100: Data_out <= 16'hDC8A	;
				14'b10001011011101: Data_out <= 16'hDC7E	;
				14'b10001011011110: Data_out <= 16'hDC72	;
				14'b10001011011111: Data_out <= 16'hDC66	;
				14'b10001011100000: Data_out <= 16'hDC5A	;
				14'b10001011100001: Data_out <= 16'hDC4E	;
				14'b10001011100010: Data_out <= 16'hDC42	;
				14'b10001011100011: Data_out <= 16'hDC36	;
				14'b10001011100100: Data_out <= 16'hDC2A	;
				14'b10001011100101: Data_out <= 16'hDC1E	;
				14'b10001011100110: Data_out <= 16'hDC11	;
				14'b10001011100111: Data_out <= 16'hDC05	;
				14'b10001011101000: Data_out <= 16'hDBF9	;
				14'b10001011101001: Data_out <= 16'hDBED	;
				14'b10001011101010: Data_out <= 16'hDBE1	;
				14'b10001011101011: Data_out <= 16'hDBD5	;
				14'b10001011101100: Data_out <= 16'hDBC9	;
				14'b10001011101101: Data_out <= 16'hDBBD	;
				14'b10001011101110: Data_out <= 16'hDBB1	;
				14'b10001011101111: Data_out <= 16'hDBA5	;
				14'b10001011110000: Data_out <= 16'hDB99	;
				14'b10001011110001: Data_out <= 16'hDB8D	;
				14'b10001011110010: Data_out <= 16'hDB81	;
				14'b10001011110011: Data_out <= 16'hDB75	;
				14'b10001011110100: Data_out <= 16'hDB69	;
				14'b10001011110101: Data_out <= 16'hDB5D	;
				14'b10001011110110: Data_out <= 16'hDB51	;
				14'b10001011110111: Data_out <= 16'hDB45	;
				14'b10001011111000: Data_out <= 16'hDB39	;
				14'b10001011111001: Data_out <= 16'hDB2D	;
				14'b10001011111010: Data_out <= 16'hDB21	;
				14'b10001011111011: Data_out <= 16'hDB14	;
				14'b10001011111100: Data_out <= 16'hDB08	;
				14'b10001011111101: Data_out <= 16'hDAFC	;
				14'b10001011111110: Data_out <= 16'hDAF0	;
				14'b10001011111111: Data_out <= 16'hDAE4	;
				14'b10001100000000: Data_out <= 16'hDAD8	;
				14'b10001100000001: Data_out <= 16'hDACC	;
				14'b10001100000010: Data_out <= 16'hDAC0	;
				14'b10001100000011: Data_out <= 16'hDAB4	;
				14'b10001100000100: Data_out <= 16'hDAA8	;
				14'b10001100000101: Data_out <= 16'hDA9C	;
				14'b10001100000110: Data_out <= 16'hDA90	;
				14'b10001100000111: Data_out <= 16'hDA84	;
				14'b10001100001000: Data_out <= 16'hDA78	;
				14'b10001100001001: Data_out <= 16'hDA6C	;
				14'b10001100001010: Data_out <= 16'hDA60	;
				14'b10001100001011: Data_out <= 16'hDA54	;
				14'b10001100001100: Data_out <= 16'hDA48	;
				14'b10001100001101: Data_out <= 16'hDA3C	;
				14'b10001100001110: Data_out <= 16'hDA30	;
				14'b10001100001111: Data_out <= 16'hDA24	;
				14'b10001100010000: Data_out <= 16'hDA18	;
				14'b10001100010001: Data_out <= 16'hDA0C	;
				14'b10001100010010: Data_out <= 16'hDA00	;
				14'b10001100010011: Data_out <= 16'hD9F4	;
				14'b10001100010100: Data_out <= 16'hD9E8	;
				14'b10001100010101: Data_out <= 16'hD9DC	;
				14'b10001100010110: Data_out <= 16'hD9D0	;
				14'b10001100010111: Data_out <= 16'hD9C4	;
				14'b10001100011000: Data_out <= 16'hD9B8	;
				14'b10001100011001: Data_out <= 16'hD9AC	;
				14'b10001100011010: Data_out <= 16'hD9A0	;
				14'b10001100011011: Data_out <= 16'hD994	;
				14'b10001100011100: Data_out <= 16'hD988	;
				14'b10001100011101: Data_out <= 16'hD97C	;
				14'b10001100011110: Data_out <= 16'hD970	;
				14'b10001100011111: Data_out <= 16'hD964	;
				14'b10001100100000: Data_out <= 16'hD958	;
				14'b10001100100001: Data_out <= 16'hD94C	;
				14'b10001100100010: Data_out <= 16'hD940	;
				14'b10001100100011: Data_out <= 16'hD934	;
				14'b10001100100100: Data_out <= 16'hD928	;
				14'b10001100100101: Data_out <= 16'hD91C	;
				14'b10001100100110: Data_out <= 16'hD910	;
				14'b10001100100111: Data_out <= 16'hD904	;
				14'b10001100101000: Data_out <= 16'hD8F8	;
				14'b10001100101001: Data_out <= 16'hD8ED	;
				14'b10001100101010: Data_out <= 16'hD8E1	;
				14'b10001100101011: Data_out <= 16'hD8D5	;
				14'b10001100101100: Data_out <= 16'hD8C9	;
				14'b10001100101101: Data_out <= 16'hD8BD	;
				14'b10001100101110: Data_out <= 16'hD8B1	;
				14'b10001100101111: Data_out <= 16'hD8A5	;
				14'b10001100110000: Data_out <= 16'hD899	;
				14'b10001100110001: Data_out <= 16'hD88D	;
				14'b10001100110010: Data_out <= 16'hD881	;
				14'b10001100110011: Data_out <= 16'hD875	;
				14'b10001100110100: Data_out <= 16'hD869	;
				14'b10001100110101: Data_out <= 16'hD85D	;
				14'b10001100110110: Data_out <= 16'hD851	;
				14'b10001100110111: Data_out <= 16'hD845	;
				14'b10001100111000: Data_out <= 16'hD839	;
				14'b10001100111001: Data_out <= 16'hD82D	;
				14'b10001100111010: Data_out <= 16'hD821	;
				14'b10001100111011: Data_out <= 16'hD815	;
				14'b10001100111100: Data_out <= 16'hD809	;
				14'b10001100111101: Data_out <= 16'hD7FD	;
				14'b10001100111110: Data_out <= 16'hD7F2	;
				14'b10001100111111: Data_out <= 16'hD7E6	;
				14'b10001101000000: Data_out <= 16'hD7DA	;
				14'b10001101000001: Data_out <= 16'hD7CE	;
				14'b10001101000010: Data_out <= 16'hD7C2	;
				14'b10001101000011: Data_out <= 16'hD7B6	;
				14'b10001101000100: Data_out <= 16'hD7AA	;
				14'b10001101000101: Data_out <= 16'hD79E	;
				14'b10001101000110: Data_out <= 16'hD792	;
				14'b10001101000111: Data_out <= 16'hD786	;
				14'b10001101001000: Data_out <= 16'hD77A	;
				14'b10001101001001: Data_out <= 16'hD76E	;
				14'b10001101001010: Data_out <= 16'hD762	;
				14'b10001101001011: Data_out <= 16'hD757	;
				14'b10001101001100: Data_out <= 16'hD74B	;
				14'b10001101001101: Data_out <= 16'hD73F	;
				14'b10001101001110: Data_out <= 16'hD733	;
				14'b10001101001111: Data_out <= 16'hD727	;
				14'b10001101010000: Data_out <= 16'hD71B	;
				14'b10001101010001: Data_out <= 16'hD70F	;
				14'b10001101010010: Data_out <= 16'hD703	;
				14'b10001101010011: Data_out <= 16'hD6F7	;
				14'b10001101010100: Data_out <= 16'hD6EB	;
				14'b10001101010101: Data_out <= 16'hD6DF	;
				14'b10001101010110: Data_out <= 16'hD6D4	;
				14'b10001101010111: Data_out <= 16'hD6C8	;
				14'b10001101011000: Data_out <= 16'hD6BC	;
				14'b10001101011001: Data_out <= 16'hD6B0	;
				14'b10001101011010: Data_out <= 16'hD6A4	;
				14'b10001101011011: Data_out <= 16'hD698	;
				14'b10001101011100: Data_out <= 16'hD68C	;
				14'b10001101011101: Data_out <= 16'hD680	;
				14'b10001101011110: Data_out <= 16'hD674	;
				14'b10001101011111: Data_out <= 16'hD669	;
				14'b10001101100000: Data_out <= 16'hD65D	;
				14'b10001101100001: Data_out <= 16'hD651	;
				14'b10001101100010: Data_out <= 16'hD645	;
				14'b10001101100011: Data_out <= 16'hD639	;
				14'b10001101100100: Data_out <= 16'hD62D	;
				14'b10001101100101: Data_out <= 16'hD621	;
				14'b10001101100110: Data_out <= 16'hD615	;
				14'b10001101100111: Data_out <= 16'hD60A	;
				14'b10001101101000: Data_out <= 16'hD5FE	;
				14'b10001101101001: Data_out <= 16'hD5F2	;
				14'b10001101101010: Data_out <= 16'hD5E6	;
				14'b10001101101011: Data_out <= 16'hD5DA	;
				14'b10001101101100: Data_out <= 16'hD5CE	;
				14'b10001101101101: Data_out <= 16'hD5C2	;
				14'b10001101101110: Data_out <= 16'hD5B6	;
				14'b10001101101111: Data_out <= 16'hD5AB	;
				14'b10001101110000: Data_out <= 16'hD59F	;
				14'b10001101110001: Data_out <= 16'hD593	;
				14'b10001101110010: Data_out <= 16'hD587	;
				14'b10001101110011: Data_out <= 16'hD57B	;
				14'b10001101110100: Data_out <= 16'hD56F	;
				14'b10001101110101: Data_out <= 16'hD563	;
				14'b10001101110110: Data_out <= 16'hD558	;
				14'b10001101110111: Data_out <= 16'hD54C	;
				14'b10001101111000: Data_out <= 16'hD540	;
				14'b10001101111001: Data_out <= 16'hD534	;
				14'b10001101111010: Data_out <= 16'hD528	;
				14'b10001101111011: Data_out <= 16'hD51C	;
				14'b10001101111100: Data_out <= 16'hD511	;
				14'b10001101111101: Data_out <= 16'hD505	;
				14'b10001101111110: Data_out <= 16'hD4F9	;
				14'b10001101111111: Data_out <= 16'hD4ED	;
				14'b10001110000000: Data_out <= 16'hD4E1	;
				14'b10001110000001: Data_out <= 16'hD4D5	;
				14'b10001110000010: Data_out <= 16'hD4CA	;
				14'b10001110000011: Data_out <= 16'hD4BE	;
				14'b10001110000100: Data_out <= 16'hD4B2	;
				14'b10001110000101: Data_out <= 16'hD4A6	;
				14'b10001110000110: Data_out <= 16'hD49A	;
				14'b10001110000111: Data_out <= 16'hD48E	;
				14'b10001110001000: Data_out <= 16'hD483	;
				14'b10001110001001: Data_out <= 16'hD477	;
				14'b10001110001010: Data_out <= 16'hD46B	;
				14'b10001110001011: Data_out <= 16'hD45F	;
				14'b10001110001100: Data_out <= 16'hD453	;
				14'b10001110001101: Data_out <= 16'hD448	;
				14'b10001110001110: Data_out <= 16'hD43C	;
				14'b10001110001111: Data_out <= 16'hD430	;
				14'b10001110010000: Data_out <= 16'hD424	;
				14'b10001110010001: Data_out <= 16'hD418	;
				14'b10001110010010: Data_out <= 16'hD40D	;
				14'b10001110010011: Data_out <= 16'hD401	;
				14'b10001110010100: Data_out <= 16'hD3F5	;
				14'b10001110010101: Data_out <= 16'hD3E9	;
				14'b10001110010110: Data_out <= 16'hD3DD	;
				14'b10001110010111: Data_out <= 16'hD3D2	;
				14'b10001110011000: Data_out <= 16'hD3C6	;
				14'b10001110011001: Data_out <= 16'hD3BA	;
				14'b10001110011010: Data_out <= 16'hD3AE	;
				14'b10001110011011: Data_out <= 16'hD3A2	;
				14'b10001110011100: Data_out <= 16'hD397	;
				14'b10001110011101: Data_out <= 16'hD38B	;
				14'b10001110011110: Data_out <= 16'hD37F	;
				14'b10001110011111: Data_out <= 16'hD373	;
				14'b10001110100000: Data_out <= 16'hD367	;
				14'b10001110100001: Data_out <= 16'hD35C	;
				14'b10001110100010: Data_out <= 16'hD350	;
				14'b10001110100011: Data_out <= 16'hD344	;
				14'b10001110100100: Data_out <= 16'hD338	;
				14'b10001110100101: Data_out <= 16'hD32D	;
				14'b10001110100110: Data_out <= 16'hD321	;
				14'b10001110100111: Data_out <= 16'hD315	;
				14'b10001110101000: Data_out <= 16'hD309	;
				14'b10001110101001: Data_out <= 16'hD2FE	;
				14'b10001110101010: Data_out <= 16'hD2F2	;
				14'b10001110101011: Data_out <= 16'hD2E6	;
				14'b10001110101100: Data_out <= 16'hD2DA	;
				14'b10001110101101: Data_out <= 16'hD2CE	;
				14'b10001110101110: Data_out <= 16'hD2C3	;
				14'b10001110101111: Data_out <= 16'hD2B7	;
				14'b10001110110000: Data_out <= 16'hD2AB	;
				14'b10001110110001: Data_out <= 16'hD29F	;
				14'b10001110110010: Data_out <= 16'hD294	;
				14'b10001110110011: Data_out <= 16'hD288	;
				14'b10001110110100: Data_out <= 16'hD27C	;
				14'b10001110110101: Data_out <= 16'hD270	;
				14'b10001110110110: Data_out <= 16'hD265	;
				14'b10001110110111: Data_out <= 16'hD259	;
				14'b10001110111000: Data_out <= 16'hD24D	;
				14'b10001110111001: Data_out <= 16'hD242	;
				14'b10001110111010: Data_out <= 16'hD236	;
				14'b10001110111011: Data_out <= 16'hD22A	;
				14'b10001110111100: Data_out <= 16'hD21E	;
				14'b10001110111101: Data_out <= 16'hD213	;
				14'b10001110111110: Data_out <= 16'hD207	;
				14'b10001110111111: Data_out <= 16'hD1FB	;
				14'b10001111000000: Data_out <= 16'hD1EF	;
				14'b10001111000001: Data_out <= 16'hD1E4	;
				14'b10001111000010: Data_out <= 16'hD1D8	;
				14'b10001111000011: Data_out <= 16'hD1CC	;
				14'b10001111000100: Data_out <= 16'hD1C1	;
				14'b10001111000101: Data_out <= 16'hD1B5	;
				14'b10001111000110: Data_out <= 16'hD1A9	;
				14'b10001111000111: Data_out <= 16'hD19D	;
				14'b10001111001000: Data_out <= 16'hD192	;
				14'b10001111001001: Data_out <= 16'hD186	;
				14'b10001111001010: Data_out <= 16'hD17A	;
				14'b10001111001011: Data_out <= 16'hD16F	;
				14'b10001111001100: Data_out <= 16'hD163	;
				14'b10001111001101: Data_out <= 16'hD157	;
				14'b10001111001110: Data_out <= 16'hD14B	;
				14'b10001111001111: Data_out <= 16'hD140	;
				14'b10001111010000: Data_out <= 16'hD134	;
				14'b10001111010001: Data_out <= 16'hD128	;
				14'b10001111010010: Data_out <= 16'hD11D	;
				14'b10001111010011: Data_out <= 16'hD111	;
				14'b10001111010100: Data_out <= 16'hD105	;
				14'b10001111010101: Data_out <= 16'hD0FA	;
				14'b10001111010110: Data_out <= 16'hD0EE	;
				14'b10001111010111: Data_out <= 16'hD0E2	;
				14'b10001111011000: Data_out <= 16'hD0D7	;
				14'b10001111011001: Data_out <= 16'hD0CB	;
				14'b10001111011010: Data_out <= 16'hD0BF	;
				14'b10001111011011: Data_out <= 16'hD0B4	;
				14'b10001111011100: Data_out <= 16'hD0A8	;
				14'b10001111011101: Data_out <= 16'hD09C	;
				14'b10001111011110: Data_out <= 16'hD090	;
				14'b10001111011111: Data_out <= 16'hD085	;
				14'b10001111100000: Data_out <= 16'hD079	;
				14'b10001111100001: Data_out <= 16'hD06D	;
				14'b10001111100010: Data_out <= 16'hD062	;
				14'b10001111100011: Data_out <= 16'hD056	;
				14'b10001111100100: Data_out <= 16'hD04A	;
				14'b10001111100101: Data_out <= 16'hD03F	;
				14'b10001111100110: Data_out <= 16'hD033	;
				14'b10001111100111: Data_out <= 16'hD028	;
				14'b10001111101000: Data_out <= 16'hD01C	;
				14'b10001111101001: Data_out <= 16'hD010	;
				14'b10001111101010: Data_out <= 16'hD005	;
				14'b10001111101011: Data_out <= 16'hCFF9	;
				14'b10001111101100: Data_out <= 16'hCFED	;
				14'b10001111101101: Data_out <= 16'hCFE2	;
				14'b10001111101110: Data_out <= 16'hCFD6	;
				14'b10001111101111: Data_out <= 16'hCFCA	;
				14'b10001111110000: Data_out <= 16'hCFBF	;
				14'b10001111110001: Data_out <= 16'hCFB3	;
				14'b10001111110010: Data_out <= 16'hCFA7	;
				14'b10001111110011: Data_out <= 16'hCF9C	;
				14'b10001111110100: Data_out <= 16'hCF90	;
				14'b10001111110101: Data_out <= 16'hCF85	;
				14'b10001111110110: Data_out <= 16'hCF79	;
				14'b10001111110111: Data_out <= 16'hCF6D	;
				14'b10001111111000: Data_out <= 16'hCF62	;
				14'b10001111111001: Data_out <= 16'hCF56	;
				14'b10001111111010: Data_out <= 16'hCF4A	;
				14'b10001111111011: Data_out <= 16'hCF3F	;
				14'b10001111111100: Data_out <= 16'hCF33	;
				14'b10001111111101: Data_out <= 16'hCF28	;
				14'b10001111111110: Data_out <= 16'hCF1C	;
				14'b10001111111111: Data_out <= 16'hCF10	;
				14'b10010000000000: Data_out <= 16'hCF05	;
				14'b10010000000001: Data_out <= 16'hCEF9	;
				14'b10010000000010: Data_out <= 16'hCEED	;
				14'b10010000000011: Data_out <= 16'hCEE2	;
				14'b10010000000100: Data_out <= 16'hCED6	;
				14'b10010000000101: Data_out <= 16'hCECB	;
				14'b10010000000110: Data_out <= 16'hCEBF	;
				14'b10010000000111: Data_out <= 16'hCEB3	;
				14'b10010000001000: Data_out <= 16'hCEA8	;
				14'b10010000001001: Data_out <= 16'hCE9C	;
				14'b10010000001010: Data_out <= 16'hCE91	;
				14'b10010000001011: Data_out <= 16'hCE85	;
				14'b10010000001100: Data_out <= 16'hCE7A	;
				14'b10010000001101: Data_out <= 16'hCE6E	;
				14'b10010000001110: Data_out <= 16'hCE62	;
				14'b10010000001111: Data_out <= 16'hCE57	;
				14'b10010000010000: Data_out <= 16'hCE4B	;
				14'b10010000010001: Data_out <= 16'hCE40	;
				14'b10010000010010: Data_out <= 16'hCE34	;
				14'b10010000010011: Data_out <= 16'hCE28	;
				14'b10010000010100: Data_out <= 16'hCE1D	;
				14'b10010000010101: Data_out <= 16'hCE11	;
				14'b10010000010110: Data_out <= 16'hCE06	;
				14'b10010000010111: Data_out <= 16'hCDFA	;
				14'b10010000011000: Data_out <= 16'hCDEF	;
				14'b10010000011001: Data_out <= 16'hCDE3	;
				14'b10010000011010: Data_out <= 16'hCDD7	;
				14'b10010000011011: Data_out <= 16'hCDCC	;
				14'b10010000011100: Data_out <= 16'hCDC0	;
				14'b10010000011101: Data_out <= 16'hCDB5	;
				14'b10010000011110: Data_out <= 16'hCDA9	;
				14'b10010000011111: Data_out <= 16'hCD9E	;
				14'b10010000100000: Data_out <= 16'hCD92	;
				14'b10010000100001: Data_out <= 16'hCD87	;
				14'b10010000100010: Data_out <= 16'hCD7B	;
				14'b10010000100011: Data_out <= 16'hCD70	;
				14'b10010000100100: Data_out <= 16'hCD64	;
				14'b10010000100101: Data_out <= 16'hCD58	;
				14'b10010000100110: Data_out <= 16'hCD4D	;
				14'b10010000100111: Data_out <= 16'hCD41	;
				14'b10010000101000: Data_out <= 16'hCD36	;
				14'b10010000101001: Data_out <= 16'hCD2A	;
				14'b10010000101010: Data_out <= 16'hCD1F	;
				14'b10010000101011: Data_out <= 16'hCD13	;
				14'b10010000101100: Data_out <= 16'hCD08	;
				14'b10010000101101: Data_out <= 16'hCCFC	;
				14'b10010000101110: Data_out <= 16'hCCF1	;
				14'b10010000101111: Data_out <= 16'hCCE5	;
				14'b10010000110000: Data_out <= 16'hCCDA	;
				14'b10010000110001: Data_out <= 16'hCCCE	;
				14'b10010000110010: Data_out <= 16'hCCC3	;
				14'b10010000110011: Data_out <= 16'hCCB7	;
				14'b10010000110100: Data_out <= 16'hCCAC	;
				14'b10010000110101: Data_out <= 16'hCCA0	;
				14'b10010000110110: Data_out <= 16'hCC95	;
				14'b10010000110111: Data_out <= 16'hCC89	;
				14'b10010000111000: Data_out <= 16'hCC7E	;
				14'b10010000111001: Data_out <= 16'hCC72	;
				14'b10010000111010: Data_out <= 16'hCC67	;
				14'b10010000111011: Data_out <= 16'hCC5B	;
				14'b10010000111100: Data_out <= 16'hCC50	;
				14'b10010000111101: Data_out <= 16'hCC44	;
				14'b10010000111110: Data_out <= 16'hCC39	;
				14'b10010000111111: Data_out <= 16'hCC2D	;
				14'b10010001000000: Data_out <= 16'hCC22	;
				14'b10010001000001: Data_out <= 16'hCC16	;
				14'b10010001000010: Data_out <= 16'hCC0B	;
				14'b10010001000011: Data_out <= 16'hCBFF	;
				14'b10010001000100: Data_out <= 16'hCBF4	;
				14'b10010001000101: Data_out <= 16'hCBE8	;
				14'b10010001000110: Data_out <= 16'hCBDD	;
				14'b10010001000111: Data_out <= 16'hCBD1	;
				14'b10010001001000: Data_out <= 16'hCBC6	;
				14'b10010001001001: Data_out <= 16'hCBBA	;
				14'b10010001001010: Data_out <= 16'hCBAF	;
				14'b10010001001011: Data_out <= 16'hCBA3	;
				14'b10010001001100: Data_out <= 16'hCB98	;
				14'b10010001001101: Data_out <= 16'hCB8C	;
				14'b10010001001110: Data_out <= 16'hCB81	;
				14'b10010001001111: Data_out <= 16'hCB75	;
				14'b10010001010000: Data_out <= 16'hCB6A	;
				14'b10010001010001: Data_out <= 16'hCB5F	;
				14'b10010001010010: Data_out <= 16'hCB53	;
				14'b10010001010011: Data_out <= 16'hCB48	;
				14'b10010001010100: Data_out <= 16'hCB3C	;
				14'b10010001010101: Data_out <= 16'hCB31	;
				14'b10010001010110: Data_out <= 16'hCB25	;
				14'b10010001010111: Data_out <= 16'hCB1A	;
				14'b10010001011000: Data_out <= 16'hCB0E	;
				14'b10010001011001: Data_out <= 16'hCB03	;
				14'b10010001011010: Data_out <= 16'hCAF8	;
				14'b10010001011011: Data_out <= 16'hCAEC	;
				14'b10010001011100: Data_out <= 16'hCAE1	;
				14'b10010001011101: Data_out <= 16'hCAD5	;
				14'b10010001011110: Data_out <= 16'hCACA	;
				14'b10010001011111: Data_out <= 16'hCABE	;
				14'b10010001100000: Data_out <= 16'hCAB3	;
				14'b10010001100001: Data_out <= 16'hCAA8	;
				14'b10010001100010: Data_out <= 16'hCA9C	;
				14'b10010001100011: Data_out <= 16'hCA91	;
				14'b10010001100100: Data_out <= 16'hCA85	;
				14'b10010001100101: Data_out <= 16'hCA7A	;
				14'b10010001100110: Data_out <= 16'hCA6E	;
				14'b10010001100111: Data_out <= 16'hCA63	;
				14'b10010001101000: Data_out <= 16'hCA58	;
				14'b10010001101001: Data_out <= 16'hCA4C	;
				14'b10010001101010: Data_out <= 16'hCA41	;
				14'b10010001101011: Data_out <= 16'hCA35	;
				14'b10010001101100: Data_out <= 16'hCA2A	;
				14'b10010001101101: Data_out <= 16'hCA1F	;
				14'b10010001101110: Data_out <= 16'hCA13	;
				14'b10010001101111: Data_out <= 16'hCA08	;
				14'b10010001110000: Data_out <= 16'hC9FC	;
				14'b10010001110001: Data_out <= 16'hC9F1	;
				14'b10010001110010: Data_out <= 16'hC9E6	;
				14'b10010001110011: Data_out <= 16'hC9DA	;
				14'b10010001110100: Data_out <= 16'hC9CF	;
				14'b10010001110101: Data_out <= 16'hC9C3	;
				14'b10010001110110: Data_out <= 16'hC9B8	;
				14'b10010001110111: Data_out <= 16'hC9AD	;
				14'b10010001111000: Data_out <= 16'hC9A1	;
				14'b10010001111001: Data_out <= 16'hC996	;
				14'b10010001111010: Data_out <= 16'hC98B	;
				14'b10010001111011: Data_out <= 16'hC97F	;
				14'b10010001111100: Data_out <= 16'hC974	;
				14'b10010001111101: Data_out <= 16'hC968	;
				14'b10010001111110: Data_out <= 16'hC95D	;
				14'b10010001111111: Data_out <= 16'hC952	;
				14'b10010010000000: Data_out <= 16'hC946	;
				14'b10010010000001: Data_out <= 16'hC93B	;
				14'b10010010000010: Data_out <= 16'hC930	;
				14'b10010010000011: Data_out <= 16'hC924	;
				14'b10010010000100: Data_out <= 16'hC919	;
				14'b10010010000101: Data_out <= 16'hC90E	;
				14'b10010010000110: Data_out <= 16'hC902	;
				14'b10010010000111: Data_out <= 16'hC8F7	;
				14'b10010010001000: Data_out <= 16'hC8EC	;
				14'b10010010001001: Data_out <= 16'hC8E0	;
				14'b10010010001010: Data_out <= 16'hC8D5	;
				14'b10010010001011: Data_out <= 16'hC8CA	;
				14'b10010010001100: Data_out <= 16'hC8BE	;
				14'b10010010001101: Data_out <= 16'hC8B3	;
				14'b10010010001110: Data_out <= 16'hC8A8	;
				14'b10010010001111: Data_out <= 16'hC89C	;
				14'b10010010010000: Data_out <= 16'hC891	;
				14'b10010010010001: Data_out <= 16'hC886	;
				14'b10010010010010: Data_out <= 16'hC87A	;
				14'b10010010010011: Data_out <= 16'hC86F	;
				14'b10010010010100: Data_out <= 16'hC864	;
				14'b10010010010101: Data_out <= 16'hC858	;
				14'b10010010010110: Data_out <= 16'hC84D	;
				14'b10010010010111: Data_out <= 16'hC842	;
				14'b10010010011000: Data_out <= 16'hC836	;
				14'b10010010011001: Data_out <= 16'hC82B	;
				14'b10010010011010: Data_out <= 16'hC820	;
				14'b10010010011011: Data_out <= 16'hC814	;
				14'b10010010011100: Data_out <= 16'hC809	;
				14'b10010010011101: Data_out <= 16'hC7FE	;
				14'b10010010011110: Data_out <= 16'hC7F3	;
				14'b10010010011111: Data_out <= 16'hC7E7	;
				14'b10010010100000: Data_out <= 16'hC7DC	;
				14'b10010010100001: Data_out <= 16'hC7D1	;
				14'b10010010100010: Data_out <= 16'hC7C5	;
				14'b10010010100011: Data_out <= 16'hC7BA	;
				14'b10010010100100: Data_out <= 16'hC7AF	;
				14'b10010010100101: Data_out <= 16'hC7A4	;
				14'b10010010100110: Data_out <= 16'hC798	;
				14'b10010010100111: Data_out <= 16'hC78D	;
				14'b10010010101000: Data_out <= 16'hC782	;
				14'b10010010101001: Data_out <= 16'hC776	;
				14'b10010010101010: Data_out <= 16'hC76B	;
				14'b10010010101011: Data_out <= 16'hC760	;
				14'b10010010101100: Data_out <= 16'hC755	;
				14'b10010010101101: Data_out <= 16'hC749	;
				14'b10010010101110: Data_out <= 16'hC73E	;
				14'b10010010101111: Data_out <= 16'hC733	;
				14'b10010010110000: Data_out <= 16'hC728	;
				14'b10010010110001: Data_out <= 16'hC71C	;
				14'b10010010110010: Data_out <= 16'hC711	;
				14'b10010010110011: Data_out <= 16'hC706	;
				14'b10010010110100: Data_out <= 16'hC6FB	;
				14'b10010010110101: Data_out <= 16'hC6EF	;
				14'b10010010110110: Data_out <= 16'hC6E4	;
				14'b10010010110111: Data_out <= 16'hC6D9	;
				14'b10010010111000: Data_out <= 16'hC6CE	;
				14'b10010010111001: Data_out <= 16'hC6C2	;
				14'b10010010111010: Data_out <= 16'hC6B7	;
				14'b10010010111011: Data_out <= 16'hC6AC	;
				14'b10010010111100: Data_out <= 16'hC6A1	;
				14'b10010010111101: Data_out <= 16'hC695	;
				14'b10010010111110: Data_out <= 16'hC68A	;
				14'b10010010111111: Data_out <= 16'hC67F	;
				14'b10010011000000: Data_out <= 16'hC674	;
				14'b10010011000001: Data_out <= 16'hC668	;
				14'b10010011000010: Data_out <= 16'hC65D	;
				14'b10010011000011: Data_out <= 16'hC652	;
				14'b10010011000100: Data_out <= 16'hC647	;
				14'b10010011000101: Data_out <= 16'hC63C	;
				14'b10010011000110: Data_out <= 16'hC630	;
				14'b10010011000111: Data_out <= 16'hC625	;
				14'b10010011001000: Data_out <= 16'hC61A	;
				14'b10010011001001: Data_out <= 16'hC60F	;
				14'b10010011001010: Data_out <= 16'hC604	;
				14'b10010011001011: Data_out <= 16'hC5F8	;
				14'b10010011001100: Data_out <= 16'hC5ED	;
				14'b10010011001101: Data_out <= 16'hC5E2	;
				14'b10010011001110: Data_out <= 16'hC5D7	;
				14'b10010011001111: Data_out <= 16'hC5CC	;
				14'b10010011010000: Data_out <= 16'hC5C0	;
				14'b10010011010001: Data_out <= 16'hC5B5	;
				14'b10010011010010: Data_out <= 16'hC5AA	;
				14'b10010011010011: Data_out <= 16'hC59F	;
				14'b10010011010100: Data_out <= 16'hC594	;
				14'b10010011010101: Data_out <= 16'hC588	;
				14'b10010011010110: Data_out <= 16'hC57D	;
				14'b10010011010111: Data_out <= 16'hC572	;
				14'b10010011011000: Data_out <= 16'hC567	;
				14'b10010011011001: Data_out <= 16'hC55C	;
				14'b10010011011010: Data_out <= 16'hC551	;
				14'b10010011011011: Data_out <= 16'hC545	;
				14'b10010011011100: Data_out <= 16'hC53A	;
				14'b10010011011101: Data_out <= 16'hC52F	;
				14'b10010011011110: Data_out <= 16'hC524	;
				14'b10010011011111: Data_out <= 16'hC519	;
				14'b10010011100000: Data_out <= 16'hC50E	;
				14'b10010011100001: Data_out <= 16'hC502	;
				14'b10010011100010: Data_out <= 16'hC4F7	;
				14'b10010011100011: Data_out <= 16'hC4EC	;
				14'b10010011100100: Data_out <= 16'hC4E1	;
				14'b10010011100101: Data_out <= 16'hC4D6	;
				14'b10010011100110: Data_out <= 16'hC4CB	;
				14'b10010011100111: Data_out <= 16'hC4C0	;
				14'b10010011101000: Data_out <= 16'hC4B4	;
				14'b10010011101001: Data_out <= 16'hC4A9	;
				14'b10010011101010: Data_out <= 16'hC49E	;
				14'b10010011101011: Data_out <= 16'hC493	;
				14'b10010011101100: Data_out <= 16'hC488	;
				14'b10010011101101: Data_out <= 16'hC47D	;
				14'b10010011101110: Data_out <= 16'hC472	;
				14'b10010011101111: Data_out <= 16'hC467	;
				14'b10010011110000: Data_out <= 16'hC45B	;
				14'b10010011110001: Data_out <= 16'hC450	;
				14'b10010011110010: Data_out <= 16'hC445	;
				14'b10010011110011: Data_out <= 16'hC43A	;
				14'b10010011110100: Data_out <= 16'hC42F	;
				14'b10010011110101: Data_out <= 16'hC424	;
				14'b10010011110110: Data_out <= 16'hC419	;
				14'b10010011110111: Data_out <= 16'hC40E	;
				14'b10010011111000: Data_out <= 16'hC403	;
				14'b10010011111001: Data_out <= 16'hC3F7	;
				14'b10010011111010: Data_out <= 16'hC3EC	;
				14'b10010011111011: Data_out <= 16'hC3E1	;
				14'b10010011111100: Data_out <= 16'hC3D6	;
				14'b10010011111101: Data_out <= 16'hC3CB	;
				14'b10010011111110: Data_out <= 16'hC3C0	;
				14'b10010011111111: Data_out <= 16'hC3B5	;
				14'b10010100000000: Data_out <= 16'hC3AA	;
				14'b10010100000001: Data_out <= 16'hC39F	;
				14'b10010100000010: Data_out <= 16'hC394	;
				14'b10010100000011: Data_out <= 16'hC389	;
				14'b10010100000100: Data_out <= 16'hC37E	;
				14'b10010100000101: Data_out <= 16'hC372	;
				14'b10010100000110: Data_out <= 16'hC367	;
				14'b10010100000111: Data_out <= 16'hC35C	;
				14'b10010100001000: Data_out <= 16'hC351	;
				14'b10010100001001: Data_out <= 16'hC346	;
				14'b10010100001010: Data_out <= 16'hC33B	;
				14'b10010100001011: Data_out <= 16'hC330	;
				14'b10010100001100: Data_out <= 16'hC325	;
				14'b10010100001101: Data_out <= 16'hC31A	;
				14'b10010100001110: Data_out <= 16'hC30F	;
				14'b10010100001111: Data_out <= 16'hC304	;
				14'b10010100010000: Data_out <= 16'hC2F9	;
				14'b10010100010001: Data_out <= 16'hC2EE	;
				14'b10010100010010: Data_out <= 16'hC2E3	;
				14'b10010100010011: Data_out <= 16'hC2D8	;
				14'b10010100010100: Data_out <= 16'hC2CD	;
				14'b10010100010101: Data_out <= 16'hC2C2	;
				14'b10010100010110: Data_out <= 16'hC2B7	;
				14'b10010100010111: Data_out <= 16'hC2AC	;
				14'b10010100011000: Data_out <= 16'hC2A1	;
				14'b10010100011001: Data_out <= 16'hC296	;
				14'b10010100011010: Data_out <= 16'hC28A	;
				14'b10010100011011: Data_out <= 16'hC27F	;
				14'b10010100011100: Data_out <= 16'hC274	;
				14'b10010100011101: Data_out <= 16'hC269	;
				14'b10010100011110: Data_out <= 16'hC25E	;
				14'b10010100011111: Data_out <= 16'hC253	;
				14'b10010100100000: Data_out <= 16'hC248	;
				14'b10010100100001: Data_out <= 16'hC23D	;
				14'b10010100100010: Data_out <= 16'hC232	;
				14'b10010100100011: Data_out <= 16'hC227	;
				14'b10010100100100: Data_out <= 16'hC21C	;
				14'b10010100100101: Data_out <= 16'hC211	;
				14'b10010100100110: Data_out <= 16'hC206	;
				14'b10010100100111: Data_out <= 16'hC1FB	;
				14'b10010100101000: Data_out <= 16'hC1F0	;
				14'b10010100101001: Data_out <= 16'hC1E5	;
				14'b10010100101010: Data_out <= 16'hC1DA	;
				14'b10010100101011: Data_out <= 16'hC1CF	;
				14'b10010100101100: Data_out <= 16'hC1C4	;
				14'b10010100101101: Data_out <= 16'hC1B9	;
				14'b10010100101110: Data_out <= 16'hC1AE	;
				14'b10010100101111: Data_out <= 16'hC1A4	;
				14'b10010100110000: Data_out <= 16'hC199	;
				14'b10010100110001: Data_out <= 16'hC18E	;
				14'b10010100110010: Data_out <= 16'hC183	;
				14'b10010100110011: Data_out <= 16'hC178	;
				14'b10010100110100: Data_out <= 16'hC16D	;
				14'b10010100110101: Data_out <= 16'hC162	;
				14'b10010100110110: Data_out <= 16'hC157	;
				14'b10010100110111: Data_out <= 16'hC14C	;
				14'b10010100111000: Data_out <= 16'hC141	;
				14'b10010100111001: Data_out <= 16'hC136	;
				14'b10010100111010: Data_out <= 16'hC12B	;
				14'b10010100111011: Data_out <= 16'hC120	;
				14'b10010100111100: Data_out <= 16'hC115	;
				14'b10010100111101: Data_out <= 16'hC10A	;
				14'b10010100111110: Data_out <= 16'hC0FF	;
				14'b10010100111111: Data_out <= 16'hC0F4	;
				14'b10010101000000: Data_out <= 16'hC0E9	;
				14'b10010101000001: Data_out <= 16'hC0DE	;
				14'b10010101000010: Data_out <= 16'hC0D3	;
				14'b10010101000011: Data_out <= 16'hC0C9	;
				14'b10010101000100: Data_out <= 16'hC0BE	;
				14'b10010101000101: Data_out <= 16'hC0B3	;
				14'b10010101000110: Data_out <= 16'hC0A8	;
				14'b10010101000111: Data_out <= 16'hC09D	;
				14'b10010101001000: Data_out <= 16'hC092	;
				14'b10010101001001: Data_out <= 16'hC087	;
				14'b10010101001010: Data_out <= 16'hC07C	;
				14'b10010101001011: Data_out <= 16'hC071	;
				14'b10010101001100: Data_out <= 16'hC066	;
				14'b10010101001101: Data_out <= 16'hC05B	;
				14'b10010101001110: Data_out <= 16'hC050	;
				14'b10010101001111: Data_out <= 16'hC046	;
				14'b10010101010000: Data_out <= 16'hC03B	;
				14'b10010101010001: Data_out <= 16'hC030	;
				14'b10010101010010: Data_out <= 16'hC025	;
				14'b10010101010011: Data_out <= 16'hC01A	;
				14'b10010101010100: Data_out <= 16'hC00F	;
				14'b10010101010101: Data_out <= 16'hC004	;
				14'b10010101010110: Data_out <= 16'hBFF9	;
				14'b10010101010111: Data_out <= 16'hBFEE	;
				14'b10010101011000: Data_out <= 16'hBFE4	;
				14'b10010101011001: Data_out <= 16'hBFD9	;
				14'b10010101011010: Data_out <= 16'hBFCE	;
				14'b10010101011011: Data_out <= 16'hBFC3	;
				14'b10010101011100: Data_out <= 16'hBFB8	;
				14'b10010101011101: Data_out <= 16'hBFAD	;
				14'b10010101011110: Data_out <= 16'hBFA2	;
				14'b10010101011111: Data_out <= 16'hBF98	;
				14'b10010101100000: Data_out <= 16'hBF8D	;
				14'b10010101100001: Data_out <= 16'hBF82	;
				14'b10010101100010: Data_out <= 16'hBF77	;
				14'b10010101100011: Data_out <= 16'hBF6C	;
				14'b10010101100100: Data_out <= 16'hBF61	;
				14'b10010101100101: Data_out <= 16'hBF56	;
				14'b10010101100110: Data_out <= 16'hBF4C	;
				14'b10010101100111: Data_out <= 16'hBF41	;
				14'b10010101101000: Data_out <= 16'hBF36	;
				14'b10010101101001: Data_out <= 16'hBF2B	;
				14'b10010101101010: Data_out <= 16'hBF20	;
				14'b10010101101011: Data_out <= 16'hBF15	;
				14'b10010101101100: Data_out <= 16'hBF0B	;
				14'b10010101101101: Data_out <= 16'hBF00	;
				14'b10010101101110: Data_out <= 16'hBEF5	;
				14'b10010101101111: Data_out <= 16'hBEEA	;
				14'b10010101110000: Data_out <= 16'hBEDF	;
				14'b10010101110001: Data_out <= 16'hBED4	;
				14'b10010101110010: Data_out <= 16'hBECA	;
				14'b10010101110011: Data_out <= 16'hBEBF	;
				14'b10010101110100: Data_out <= 16'hBEB4	;
				14'b10010101110101: Data_out <= 16'hBEA9	;
				14'b10010101110110: Data_out <= 16'hBE9E	;
				14'b10010101110111: Data_out <= 16'hBE94	;
				14'b10010101111000: Data_out <= 16'hBE89	;
				14'b10010101111001: Data_out <= 16'hBE7E	;
				14'b10010101111010: Data_out <= 16'hBE73	;
				14'b10010101111011: Data_out <= 16'hBE68	;
				14'b10010101111100: Data_out <= 16'hBE5E	;
				14'b10010101111101: Data_out <= 16'hBE53	;
				14'b10010101111110: Data_out <= 16'hBE48	;
				14'b10010101111111: Data_out <= 16'hBE3D	;
				14'b10010110000000: Data_out <= 16'hBE32	;
				14'b10010110000001: Data_out <= 16'hBE28	;
				14'b10010110000010: Data_out <= 16'hBE1D	;
				14'b10010110000011: Data_out <= 16'hBE12	;
				14'b10010110000100: Data_out <= 16'hBE07	;
				14'b10010110000101: Data_out <= 16'hBDFD	;
				14'b10010110000110: Data_out <= 16'hBDF2	;
				14'b10010110000111: Data_out <= 16'hBDE7	;
				14'b10010110001000: Data_out <= 16'hBDDC	;
				14'b10010110001001: Data_out <= 16'hBDD2	;
				14'b10010110001010: Data_out <= 16'hBDC7	;
				14'b10010110001011: Data_out <= 16'hBDBC	;
				14'b10010110001100: Data_out <= 16'hBDB1	;
				14'b10010110001101: Data_out <= 16'hBDA7	;
				14'b10010110001110: Data_out <= 16'hBD9C	;
				14'b10010110001111: Data_out <= 16'hBD91	;
				14'b10010110010000: Data_out <= 16'hBD86	;
				14'b10010110010001: Data_out <= 16'hBD7C	;
				14'b10010110010010: Data_out <= 16'hBD71	;
				14'b10010110010011: Data_out <= 16'hBD66	;
				14'b10010110010100: Data_out <= 16'hBD5B	;
				14'b10010110010101: Data_out <= 16'hBD51	;
				14'b10010110010110: Data_out <= 16'hBD46	;
				14'b10010110010111: Data_out <= 16'hBD3B	;
				14'b10010110011000: Data_out <= 16'hBD31	;
				14'b10010110011001: Data_out <= 16'hBD26	;
				14'b10010110011010: Data_out <= 16'hBD1B	;
				14'b10010110011011: Data_out <= 16'hBD10	;
				14'b10010110011100: Data_out <= 16'hBD06	;
				14'b10010110011101: Data_out <= 16'hBCFB	;
				14'b10010110011110: Data_out <= 16'hBCF0	;
				14'b10010110011111: Data_out <= 16'hBCE6	;
				14'b10010110100000: Data_out <= 16'hBCDB	;
				14'b10010110100001: Data_out <= 16'hBCD0	;
				14'b10010110100010: Data_out <= 16'hBCC5	;
				14'b10010110100011: Data_out <= 16'hBCBB	;
				14'b10010110100100: Data_out <= 16'hBCB0	;
				14'b10010110100101: Data_out <= 16'hBCA5	;
				14'b10010110100110: Data_out <= 16'hBC9B	;
				14'b10010110100111: Data_out <= 16'hBC90	;
				14'b10010110101000: Data_out <= 16'hBC85	;
				14'b10010110101001: Data_out <= 16'hBC7B	;
				14'b10010110101010: Data_out <= 16'hBC70	;
				14'b10010110101011: Data_out <= 16'hBC65	;
				14'b10010110101100: Data_out <= 16'hBC5B	;
				14'b10010110101101: Data_out <= 16'hBC50	;
				14'b10010110101110: Data_out <= 16'hBC45	;
				14'b10010110101111: Data_out <= 16'hBC3B	;
				14'b10010110110000: Data_out <= 16'hBC30	;
				14'b10010110110001: Data_out <= 16'hBC25	;
				14'b10010110110010: Data_out <= 16'hBC1B	;
				14'b10010110110011: Data_out <= 16'hBC10	;
				14'b10010110110100: Data_out <= 16'hBC05	;
				14'b10010110110101: Data_out <= 16'hBBFB	;
				14'b10010110110110: Data_out <= 16'hBBF0	;
				14'b10010110110111: Data_out <= 16'hBBE5	;
				14'b10010110111000: Data_out <= 16'hBBDB	;
				14'b10010110111001: Data_out <= 16'hBBD0	;
				14'b10010110111010: Data_out <= 16'hBBC6	;
				14'b10010110111011: Data_out <= 16'hBBBB	;
				14'b10010110111100: Data_out <= 16'hBBB0	;
				14'b10010110111101: Data_out <= 16'hBBA6	;
				14'b10010110111110: Data_out <= 16'hBB9B	;
				14'b10010110111111: Data_out <= 16'hBB90	;
				14'b10010111000000: Data_out <= 16'hBB86	;
				14'b10010111000001: Data_out <= 16'hBB7B	;
				14'b10010111000010: Data_out <= 16'hBB71	;
				14'b10010111000011: Data_out <= 16'hBB66	;
				14'b10010111000100: Data_out <= 16'hBB5B	;
				14'b10010111000101: Data_out <= 16'hBB51	;
				14'b10010111000110: Data_out <= 16'hBB46	;
				14'b10010111000111: Data_out <= 16'hBB3C	;
				14'b10010111001000: Data_out <= 16'hBB31	;
				14'b10010111001001: Data_out <= 16'hBB26	;
				14'b10010111001010: Data_out <= 16'hBB1C	;
				14'b10010111001011: Data_out <= 16'hBB11	;
				14'b10010111001100: Data_out <= 16'hBB07	;
				14'b10010111001101: Data_out <= 16'hBAFC	;
				14'b10010111001110: Data_out <= 16'hBAF1	;
				14'b10010111001111: Data_out <= 16'hBAE7	;
				14'b10010111010000: Data_out <= 16'hBADC	;
				14'b10010111010001: Data_out <= 16'hBAD2	;
				14'b10010111010010: Data_out <= 16'hBAC7	;
				14'b10010111010011: Data_out <= 16'hBABD	;
				14'b10010111010100: Data_out <= 16'hBAB2	;
				14'b10010111010101: Data_out <= 16'hBAA7	;
				14'b10010111010110: Data_out <= 16'hBA9D	;
				14'b10010111010111: Data_out <= 16'hBA92	;
				14'b10010111011000: Data_out <= 16'hBA88	;
				14'b10010111011001: Data_out <= 16'hBA7D	;
				14'b10010111011010: Data_out <= 16'hBA73	;
				14'b10010111011011: Data_out <= 16'hBA68	;
				14'b10010111011100: Data_out <= 16'hBA5E	;
				14'b10010111011101: Data_out <= 16'hBA53	;
				14'b10010111011110: Data_out <= 16'hBA49	;
				14'b10010111011111: Data_out <= 16'hBA3E	;
				14'b10010111100000: Data_out <= 16'hBA33	;
				14'b10010111100001: Data_out <= 16'hBA29	;
				14'b10010111100010: Data_out <= 16'hBA1E	;
				14'b10010111100011: Data_out <= 16'hBA14	;
				14'b10010111100100: Data_out <= 16'hBA09	;
				14'b10010111100101: Data_out <= 16'hB9FF	;
				14'b10010111100110: Data_out <= 16'hB9F4	;
				14'b10010111100111: Data_out <= 16'hB9EA	;
				14'b10010111101000: Data_out <= 16'hB9DF	;
				14'b10010111101001: Data_out <= 16'hB9D5	;
				14'b10010111101010: Data_out <= 16'hB9CA	;
				14'b10010111101011: Data_out <= 16'hB9C0	;
				14'b10010111101100: Data_out <= 16'hB9B5	;
				14'b10010111101101: Data_out <= 16'hB9AB	;
				14'b10010111101110: Data_out <= 16'hB9A0	;
				14'b10010111101111: Data_out <= 16'hB996	;
				14'b10010111110000: Data_out <= 16'hB98B	;
				14'b10010111110001: Data_out <= 16'hB981	;
				14'b10010111110010: Data_out <= 16'hB976	;
				14'b10010111110011: Data_out <= 16'hB96C	;
				14'b10010111110100: Data_out <= 16'hB961	;
				14'b10010111110101: Data_out <= 16'hB957	;
				14'b10010111110110: Data_out <= 16'hB94C	;
				14'b10010111110111: Data_out <= 16'hB942	;
				14'b10010111111000: Data_out <= 16'hB937	;
				14'b10010111111001: Data_out <= 16'hB92D	;
				14'b10010111111010: Data_out <= 16'hB922	;
				14'b10010111111011: Data_out <= 16'hB918	;
				14'b10010111111100: Data_out <= 16'hB90E	;
				14'b10010111111101: Data_out <= 16'hB903	;
				14'b10010111111110: Data_out <= 16'hB8F9	;
				14'b10010111111111: Data_out <= 16'hB8EE	;
				14'b10011000000000: Data_out <= 16'hB8E4	;
				14'b10011000000001: Data_out <= 16'hB8D9	;
				14'b10011000000010: Data_out <= 16'hB8CF	;
				14'b10011000000011: Data_out <= 16'hB8C4	;
				14'b10011000000100: Data_out <= 16'hB8BA	;
				14'b10011000000101: Data_out <= 16'hB8B0	;
				14'b10011000000110: Data_out <= 16'hB8A5	;
				14'b10011000000111: Data_out <= 16'hB89B	;
				14'b10011000001000: Data_out <= 16'hB890	;
				14'b10011000001001: Data_out <= 16'hB886	;
				14'b10011000001010: Data_out <= 16'hB87B	;
				14'b10011000001011: Data_out <= 16'hB871	;
				14'b10011000001100: Data_out <= 16'hB867	;
				14'b10011000001101: Data_out <= 16'hB85C	;
				14'b10011000001110: Data_out <= 16'hB852	;
				14'b10011000001111: Data_out <= 16'hB847	;
				14'b10011000010000: Data_out <= 16'hB83D	;
				14'b10011000010001: Data_out <= 16'hB832	;
				14'b10011000010010: Data_out <= 16'hB828	;
				14'b10011000010011: Data_out <= 16'hB81E	;
				14'b10011000010100: Data_out <= 16'hB813	;
				14'b10011000010101: Data_out <= 16'hB809	;
				14'b10011000010110: Data_out <= 16'hB7FF	;
				14'b10011000010111: Data_out <= 16'hB7F4	;
				14'b10011000011000: Data_out <= 16'hB7EA	;
				14'b10011000011001: Data_out <= 16'hB7DF	;
				14'b10011000011010: Data_out <= 16'hB7D5	;
				14'b10011000011011: Data_out <= 16'hB7CB	;
				14'b10011000011100: Data_out <= 16'hB7C0	;
				14'b10011000011101: Data_out <= 16'hB7B6	;
				14'b10011000011110: Data_out <= 16'hB7AB	;
				14'b10011000011111: Data_out <= 16'hB7A1	;
				14'b10011000100000: Data_out <= 16'hB797	;
				14'b10011000100001: Data_out <= 16'hB78C	;
				14'b10011000100010: Data_out <= 16'hB782	;
				14'b10011000100011: Data_out <= 16'hB778	;
				14'b10011000100100: Data_out <= 16'hB76D	;
				14'b10011000100101: Data_out <= 16'hB763	;
				14'b10011000100110: Data_out <= 16'hB759	;
				14'b10011000100111: Data_out <= 16'hB74E	;
				14'b10011000101000: Data_out <= 16'hB744	;
				14'b10011000101001: Data_out <= 16'hB73A	;
				14'b10011000101010: Data_out <= 16'hB72F	;
				14'b10011000101011: Data_out <= 16'hB725	;
				14'b10011000101100: Data_out <= 16'hB71B	;
				14'b10011000101101: Data_out <= 16'hB710	;
				14'b10011000101110: Data_out <= 16'hB706	;
				14'b10011000101111: Data_out <= 16'hB6FC	;
				14'b10011000110000: Data_out <= 16'hB6F1	;
				14'b10011000110001: Data_out <= 16'hB6E7	;
				14'b10011000110010: Data_out <= 16'hB6DD	;
				14'b10011000110011: Data_out <= 16'hB6D2	;
				14'b10011000110100: Data_out <= 16'hB6C8	;
				14'b10011000110101: Data_out <= 16'hB6BE	;
				14'b10011000110110: Data_out <= 16'hB6B3	;
				14'b10011000110111: Data_out <= 16'hB6A9	;
				14'b10011000111000: Data_out <= 16'hB69F	;
				14'b10011000111001: Data_out <= 16'hB695	;
				14'b10011000111010: Data_out <= 16'hB68A	;
				14'b10011000111011: Data_out <= 16'hB680	;
				14'b10011000111100: Data_out <= 16'hB676	;
				14'b10011000111101: Data_out <= 16'hB66B	;
				14'b10011000111110: Data_out <= 16'hB661	;
				14'b10011000111111: Data_out <= 16'hB657	;
				14'b10011001000000: Data_out <= 16'hB64D	;
				14'b10011001000001: Data_out <= 16'hB642	;
				14'b10011001000010: Data_out <= 16'hB638	;
				14'b10011001000011: Data_out <= 16'hB62E	;
				14'b10011001000100: Data_out <= 16'hB624	;
				14'b10011001000101: Data_out <= 16'hB619	;
				14'b10011001000110: Data_out <= 16'hB60F	;
				14'b10011001000111: Data_out <= 16'hB605	;
				14'b10011001001000: Data_out <= 16'hB5FA	;
				14'b10011001001001: Data_out <= 16'hB5F0	;
				14'b10011001001010: Data_out <= 16'hB5E6	;
				14'b10011001001011: Data_out <= 16'hB5DC	;
				14'b10011001001100: Data_out <= 16'hB5D2	;
				14'b10011001001101: Data_out <= 16'hB5C7	;
				14'b10011001001110: Data_out <= 16'hB5BD	;
				14'b10011001001111: Data_out <= 16'hB5B3	;
				14'b10011001010000: Data_out <= 16'hB5A9	;
				14'b10011001010001: Data_out <= 16'hB59E	;
				14'b10011001010010: Data_out <= 16'hB594	;
				14'b10011001010011: Data_out <= 16'hB58A	;
				14'b10011001010100: Data_out <= 16'hB580	;
				14'b10011001010101: Data_out <= 16'hB575	;
				14'b10011001010110: Data_out <= 16'hB56B	;
				14'b10011001010111: Data_out <= 16'hB561	;
				14'b10011001011000: Data_out <= 16'hB557	;
				14'b10011001011001: Data_out <= 16'hB54D	;
				14'b10011001011010: Data_out <= 16'hB542	;
				14'b10011001011011: Data_out <= 16'hB538	;
				14'b10011001011100: Data_out <= 16'hB52E	;
				14'b10011001011101: Data_out <= 16'hB524	;
				14'b10011001011110: Data_out <= 16'hB51A	;
				14'b10011001011111: Data_out <= 16'hB50F	;
				14'b10011001100000: Data_out <= 16'hB505	;
				14'b10011001100001: Data_out <= 16'hB4FB	;
				14'b10011001100010: Data_out <= 16'hB4F1	;
				14'b10011001100011: Data_out <= 16'hB4E7	;
				14'b10011001100100: Data_out <= 16'hB4DD	;
				14'b10011001100101: Data_out <= 16'hB4D2	;
				14'b10011001100110: Data_out <= 16'hB4C8	;
				14'b10011001100111: Data_out <= 16'hB4BE	;
				14'b10011001101000: Data_out <= 16'hB4B4	;
				14'b10011001101001: Data_out <= 16'hB4AA	;
				14'b10011001101010: Data_out <= 16'hB4A0	;
				14'b10011001101011: Data_out <= 16'hB495	;
				14'b10011001101100: Data_out <= 16'hB48B	;
				14'b10011001101101: Data_out <= 16'hB481	;
				14'b10011001101110: Data_out <= 16'hB477	;
				14'b10011001101111: Data_out <= 16'hB46D	;
				14'b10011001110000: Data_out <= 16'hB463	;
				14'b10011001110001: Data_out <= 16'hB459	;
				14'b10011001110010: Data_out <= 16'hB44E	;
				14'b10011001110011: Data_out <= 16'hB444	;
				14'b10011001110100: Data_out <= 16'hB43A	;
				14'b10011001110101: Data_out <= 16'hB430	;
				14'b10011001110110: Data_out <= 16'hB426	;
				14'b10011001110111: Data_out <= 16'hB41C	;
				14'b10011001111000: Data_out <= 16'hB412	;
				14'b10011001111001: Data_out <= 16'hB408	;
				14'b10011001111010: Data_out <= 16'hB3FD	;
				14'b10011001111011: Data_out <= 16'hB3F3	;
				14'b10011001111100: Data_out <= 16'hB3E9	;
				14'b10011001111101: Data_out <= 16'hB3DF	;
				14'b10011001111110: Data_out <= 16'hB3D5	;
				14'b10011001111111: Data_out <= 16'hB3CB	;
				14'b10011010000000: Data_out <= 16'hB3C1	;
				14'b10011010000001: Data_out <= 16'hB3B7	;
				14'b10011010000010: Data_out <= 16'hB3AD	;
				14'b10011010000011: Data_out <= 16'hB3A3	;
				14'b10011010000100: Data_out <= 16'hB398	;
				14'b10011010000101: Data_out <= 16'hB38E	;
				14'b10011010000110: Data_out <= 16'hB384	;
				14'b10011010000111: Data_out <= 16'hB37A	;
				14'b10011010001000: Data_out <= 16'hB370	;
				14'b10011010001001: Data_out <= 16'hB366	;
				14'b10011010001010: Data_out <= 16'hB35C	;
				14'b10011010001011: Data_out <= 16'hB352	;
				14'b10011010001100: Data_out <= 16'hB348	;
				14'b10011010001101: Data_out <= 16'hB33E	;
				14'b10011010001110: Data_out <= 16'hB334	;
				14'b10011010001111: Data_out <= 16'hB32A	;
				14'b10011010010000: Data_out <= 16'hB320	;
				14'b10011010010001: Data_out <= 16'hB316	;
				14'b10011010010010: Data_out <= 16'hB30C	;
				14'b10011010010011: Data_out <= 16'hB302	;
				14'b10011010010100: Data_out <= 16'hB2F8	;
				14'b10011010010101: Data_out <= 16'hB2EE	;
				14'b10011010010110: Data_out <= 16'hB2E3	;
				14'b10011010010111: Data_out <= 16'hB2D9	;
				14'b10011010011000: Data_out <= 16'hB2CF	;
				14'b10011010011001: Data_out <= 16'hB2C5	;
				14'b10011010011010: Data_out <= 16'hB2BB	;
				14'b10011010011011: Data_out <= 16'hB2B1	;
				14'b10011010011100: Data_out <= 16'hB2A7	;
				14'b10011010011101: Data_out <= 16'hB29D	;
				14'b10011010011110: Data_out <= 16'hB293	;
				14'b10011010011111: Data_out <= 16'hB289	;
				14'b10011010100000: Data_out <= 16'hB27F	;
				14'b10011010100001: Data_out <= 16'hB275	;
				14'b10011010100010: Data_out <= 16'hB26B	;
				14'b10011010100011: Data_out <= 16'hB261	;
				14'b10011010100100: Data_out <= 16'hB257	;
				14'b10011010100101: Data_out <= 16'hB24D	;
				14'b10011010100110: Data_out <= 16'hB243	;
				14'b10011010100111: Data_out <= 16'hB239	;
				14'b10011010101000: Data_out <= 16'hB22F	;
				14'b10011010101001: Data_out <= 16'hB225	;
				14'b10011010101010: Data_out <= 16'hB21B	;
				14'b10011010101011: Data_out <= 16'hB211	;
				14'b10011010101100: Data_out <= 16'hB208	;
				14'b10011010101101: Data_out <= 16'hB1FE	;
				14'b10011010101110: Data_out <= 16'hB1F4	;
				14'b10011010101111: Data_out <= 16'hB1EA	;
				14'b10011010110000: Data_out <= 16'hB1E0	;
				14'b10011010110001: Data_out <= 16'hB1D6	;
				14'b10011010110010: Data_out <= 16'hB1CC	;
				14'b10011010110011: Data_out <= 16'hB1C2	;
				14'b10011010110100: Data_out <= 16'hB1B8	;
				14'b10011010110101: Data_out <= 16'hB1AE	;
				14'b10011010110110: Data_out <= 16'hB1A4	;
				14'b10011010110111: Data_out <= 16'hB19A	;
				14'b10011010111000: Data_out <= 16'hB190	;
				14'b10011010111001: Data_out <= 16'hB186	;
				14'b10011010111010: Data_out <= 16'hB17C	;
				14'b10011010111011: Data_out <= 16'hB172	;
				14'b10011010111100: Data_out <= 16'hB168	;
				14'b10011010111101: Data_out <= 16'hB15F	;
				14'b10011010111110: Data_out <= 16'hB155	;
				14'b10011010111111: Data_out <= 16'hB14B	;
				14'b10011011000000: Data_out <= 16'hB141	;
				14'b10011011000001: Data_out <= 16'hB137	;
				14'b10011011000010: Data_out <= 16'hB12D	;
				14'b10011011000011: Data_out <= 16'hB123	;
				14'b10011011000100: Data_out <= 16'hB119	;
				14'b10011011000101: Data_out <= 16'hB10F	;
				14'b10011011000110: Data_out <= 16'hB105	;
				14'b10011011000111: Data_out <= 16'hB0FC	;
				14'b10011011001000: Data_out <= 16'hB0F2	;
				14'b10011011001001: Data_out <= 16'hB0E8	;
				14'b10011011001010: Data_out <= 16'hB0DE	;
				14'b10011011001011: Data_out <= 16'hB0D4	;
				14'b10011011001100: Data_out <= 16'hB0CA	;
				14'b10011011001101: Data_out <= 16'hB0C0	;
				14'b10011011001110: Data_out <= 16'hB0B6	;
				14'b10011011001111: Data_out <= 16'hB0AD	;
				14'b10011011010000: Data_out <= 16'hB0A3	;
				14'b10011011010001: Data_out <= 16'hB099	;
				14'b10011011010010: Data_out <= 16'hB08F	;
				14'b10011011010011: Data_out <= 16'hB085	;
				14'b10011011010100: Data_out <= 16'hB07B	;
				14'b10011011010101: Data_out <= 16'hB071	;
				14'b10011011010110: Data_out <= 16'hB068	;
				14'b10011011010111: Data_out <= 16'hB05E	;
				14'b10011011011000: Data_out <= 16'hB054	;
				14'b10011011011001: Data_out <= 16'hB04A	;
				14'b10011011011010: Data_out <= 16'hB040	;
				14'b10011011011011: Data_out <= 16'hB036	;
				14'b10011011011100: Data_out <= 16'hB02D	;
				14'b10011011011101: Data_out <= 16'hB023	;
				14'b10011011011110: Data_out <= 16'hB019	;
				14'b10011011011111: Data_out <= 16'hB00F	;
				14'b10011011100000: Data_out <= 16'hB005	;
				14'b10011011100001: Data_out <= 16'hAFFC	;
				14'b10011011100010: Data_out <= 16'hAFF2	;
				14'b10011011100011: Data_out <= 16'hAFE8	;
				14'b10011011100100: Data_out <= 16'hAFDE	;
				14'b10011011100101: Data_out <= 16'hAFD4	;
				14'b10011011100110: Data_out <= 16'hAFCB	;
				14'b10011011100111: Data_out <= 16'hAFC1	;
				14'b10011011101000: Data_out <= 16'hAFB7	;
				14'b10011011101001: Data_out <= 16'hAFAD	;
				14'b10011011101010: Data_out <= 16'hAFA3	;
				14'b10011011101011: Data_out <= 16'hAF9A	;
				14'b10011011101100: Data_out <= 16'hAF90	;
				14'b10011011101101: Data_out <= 16'hAF86	;
				14'b10011011101110: Data_out <= 16'hAF7C	;
				14'b10011011101111: Data_out <= 16'hAF73	;
				14'b10011011110000: Data_out <= 16'hAF69	;
				14'b10011011110001: Data_out <= 16'hAF5F	;
				14'b10011011110010: Data_out <= 16'hAF55	;
				14'b10011011110011: Data_out <= 16'hAF4B	;
				14'b10011011110100: Data_out <= 16'hAF42	;
				14'b10011011110101: Data_out <= 16'hAF38	;
				14'b10011011110110: Data_out <= 16'hAF2E	;
				14'b10011011110111: Data_out <= 16'hAF24	;
				14'b10011011111000: Data_out <= 16'hAF1B	;
				14'b10011011111001: Data_out <= 16'hAF11	;
				14'b10011011111010: Data_out <= 16'hAF07	;
				14'b10011011111011: Data_out <= 16'hAEFE	;
				14'b10011011111100: Data_out <= 16'hAEF4	;
				14'b10011011111101: Data_out <= 16'hAEEA	;
				14'b10011011111110: Data_out <= 16'hAEE0	;
				14'b10011011111111: Data_out <= 16'hAED7	;
				14'b10011100000000: Data_out <= 16'hAECD	;
				14'b10011100000001: Data_out <= 16'hAEC3	;
				14'b10011100000010: Data_out <= 16'hAEBA	;
				14'b10011100000011: Data_out <= 16'hAEB0	;
				14'b10011100000100: Data_out <= 16'hAEA6	;
				14'b10011100000101: Data_out <= 16'hAE9C	;
				14'b10011100000110: Data_out <= 16'hAE93	;
				14'b10011100000111: Data_out <= 16'hAE89	;
				14'b10011100001000: Data_out <= 16'hAE7F	;
				14'b10011100001001: Data_out <= 16'hAE76	;
				14'b10011100001010: Data_out <= 16'hAE6C	;
				14'b10011100001011: Data_out <= 16'hAE62	;
				14'b10011100001100: Data_out <= 16'hAE59	;
				14'b10011100001101: Data_out <= 16'hAE4F	;
				14'b10011100001110: Data_out <= 16'hAE45	;
				14'b10011100001111: Data_out <= 16'hAE3C	;
				14'b10011100010000: Data_out <= 16'hAE32	;
				14'b10011100010001: Data_out <= 16'hAE28	;
				14'b10011100010010: Data_out <= 16'hAE1F	;
				14'b10011100010011: Data_out <= 16'hAE15	;
				14'b10011100010100: Data_out <= 16'hAE0B	;
				14'b10011100010101: Data_out <= 16'hAE02	;
				14'b10011100010110: Data_out <= 16'hADF8	;
				14'b10011100010111: Data_out <= 16'hADEE	;
				14'b10011100011000: Data_out <= 16'hADE5	;
				14'b10011100011001: Data_out <= 16'hADDB	;
				14'b10011100011010: Data_out <= 16'hADD1	;
				14'b10011100011011: Data_out <= 16'hADC8	;
				14'b10011100011100: Data_out <= 16'hADBE	;
				14'b10011100011101: Data_out <= 16'hADB5	;
				14'b10011100011110: Data_out <= 16'hADAB	;
				14'b10011100011111: Data_out <= 16'hADA1	;
				14'b10011100100000: Data_out <= 16'hAD98	;
				14'b10011100100001: Data_out <= 16'hAD8E	;
				14'b10011100100010: Data_out <= 16'hAD84	;
				14'b10011100100011: Data_out <= 16'hAD7B	;
				14'b10011100100100: Data_out <= 16'hAD71	;
				14'b10011100100101: Data_out <= 16'hAD68	;
				14'b10011100100110: Data_out <= 16'hAD5E	;
				14'b10011100100111: Data_out <= 16'hAD54	;
				14'b10011100101000: Data_out <= 16'hAD4B	;
				14'b10011100101001: Data_out <= 16'hAD41	;
				14'b10011100101010: Data_out <= 16'hAD38	;
				14'b10011100101011: Data_out <= 16'hAD2E	;
				14'b10011100101100: Data_out <= 16'hAD25	;
				14'b10011100101101: Data_out <= 16'hAD1B	;
				14'b10011100101110: Data_out <= 16'hAD11	;
				14'b10011100101111: Data_out <= 16'hAD08	;
				14'b10011100110000: Data_out <= 16'hACFE	;
				14'b10011100110001: Data_out <= 16'hACF5	;
				14'b10011100110010: Data_out <= 16'hACEB	;
				14'b10011100110011: Data_out <= 16'hACE2	;
				14'b10011100110100: Data_out <= 16'hACD8	;
				14'b10011100110101: Data_out <= 16'hACCE	;
				14'b10011100110110: Data_out <= 16'hACC5	;
				14'b10011100110111: Data_out <= 16'hACBB	;
				14'b10011100111000: Data_out <= 16'hACB2	;
				14'b10011100111001: Data_out <= 16'hACA8	;
				14'b10011100111010: Data_out <= 16'hAC9F	;
				14'b10011100111011: Data_out <= 16'hAC95	;
				14'b10011100111100: Data_out <= 16'hAC8C	;
				14'b10011100111101: Data_out <= 16'hAC82	;
				14'b10011100111110: Data_out <= 16'hAC79	;
				14'b10011100111111: Data_out <= 16'hAC6F	;
				14'b10011101000000: Data_out <= 16'hAC66	;
				14'b10011101000001: Data_out <= 16'hAC5C	;
				14'b10011101000010: Data_out <= 16'hAC53	;
				14'b10011101000011: Data_out <= 16'hAC49	;
				14'b10011101000100: Data_out <= 16'hAC40	;
				14'b10011101000101: Data_out <= 16'hAC36	;
				14'b10011101000110: Data_out <= 16'hAC2D	;
				14'b10011101000111: Data_out <= 16'hAC23	;
				14'b10011101001000: Data_out <= 16'hAC1A	;
				14'b10011101001001: Data_out <= 16'hAC10	;
				14'b10011101001010: Data_out <= 16'hAC07	;
				14'b10011101001011: Data_out <= 16'hABFD	;
				14'b10011101001100: Data_out <= 16'hABF4	;
				14'b10011101001101: Data_out <= 16'hABEA	;
				14'b10011101001110: Data_out <= 16'hABE1	;
				14'b10011101001111: Data_out <= 16'hABD7	;
				14'b10011101010000: Data_out <= 16'hABCE	;
				14'b10011101010001: Data_out <= 16'hABC4	;
				14'b10011101010010: Data_out <= 16'hABBB	;
				14'b10011101010011: Data_out <= 16'hABB1	;
				14'b10011101010100: Data_out <= 16'hABA8	;
				14'b10011101010101: Data_out <= 16'hAB9E	;
				14'b10011101010110: Data_out <= 16'hAB95	;
				14'b10011101010111: Data_out <= 16'hAB8C	;
				14'b10011101011000: Data_out <= 16'hAB82	;
				14'b10011101011001: Data_out <= 16'hAB79	;
				14'b10011101011010: Data_out <= 16'hAB6F	;
				14'b10011101011011: Data_out <= 16'hAB66	;
				14'b10011101011100: Data_out <= 16'hAB5C	;
				14'b10011101011101: Data_out <= 16'hAB53	;
				14'b10011101011110: Data_out <= 16'hAB4A	;
				14'b10011101011111: Data_out <= 16'hAB40	;
				14'b10011101100000: Data_out <= 16'hAB37	;
				14'b10011101100001: Data_out <= 16'hAB2D	;
				14'b10011101100010: Data_out <= 16'hAB24	;
				14'b10011101100011: Data_out <= 16'hAB1A	;
				14'b10011101100100: Data_out <= 16'hAB11	;
				14'b10011101100101: Data_out <= 16'hAB08	;
				14'b10011101100110: Data_out <= 16'hAAFE	;
				14'b10011101100111: Data_out <= 16'hAAF5	;
				14'b10011101101000: Data_out <= 16'hAAEC	;
				14'b10011101101001: Data_out <= 16'hAAE2	;
				14'b10011101101010: Data_out <= 16'hAAD9	;
				14'b10011101101011: Data_out <= 16'hAACF	;
				14'b10011101101100: Data_out <= 16'hAAC6	;
				14'b10011101101101: Data_out <= 16'hAABD	;
				14'b10011101101110: Data_out <= 16'hAAB3	;
				14'b10011101101111: Data_out <= 16'hAAAA	;
				14'b10011101110000: Data_out <= 16'hAAA1	;
				14'b10011101110001: Data_out <= 16'hAA97	;
				14'b10011101110010: Data_out <= 16'hAA8E	;
				14'b10011101110011: Data_out <= 16'hAA84	;
				14'b10011101110100: Data_out <= 16'hAA7B	;
				14'b10011101110101: Data_out <= 16'hAA72	;
				14'b10011101110110: Data_out <= 16'hAA68	;
				14'b10011101110111: Data_out <= 16'hAA5F	;
				14'b10011101111000: Data_out <= 16'hAA56	;
				14'b10011101111001: Data_out <= 16'hAA4C	;
				14'b10011101111010: Data_out <= 16'hAA43	;
				14'b10011101111011: Data_out <= 16'hAA3A	;
				14'b10011101111100: Data_out <= 16'hAA30	;
				14'b10011101111101: Data_out <= 16'hAA27	;
				14'b10011101111110: Data_out <= 16'hAA1E	;
				14'b10011101111111: Data_out <= 16'hAA14	;
				14'b10011110000000: Data_out <= 16'hAA0B	;
				14'b10011110000001: Data_out <= 16'hAA02	;
				14'b10011110000010: Data_out <= 16'hA9F9	;
				14'b10011110000011: Data_out <= 16'hA9EF	;
				14'b10011110000100: Data_out <= 16'hA9E6	;
				14'b10011110000101: Data_out <= 16'hA9DD	;
				14'b10011110000110: Data_out <= 16'hA9D3	;
				14'b10011110000111: Data_out <= 16'hA9CA	;
				14'b10011110001000: Data_out <= 16'hA9C1	;
				14'b10011110001001: Data_out <= 16'hA9B7	;
				14'b10011110001010: Data_out <= 16'hA9AE	;
				14'b10011110001011: Data_out <= 16'hA9A5	;
				14'b10011110001100: Data_out <= 16'hA99C	;
				14'b10011110001101: Data_out <= 16'hA992	;
				14'b10011110001110: Data_out <= 16'hA989	;
				14'b10011110001111: Data_out <= 16'hA980	;
				14'b10011110010000: Data_out <= 16'hA977	;
				14'b10011110010001: Data_out <= 16'hA96D	;
				14'b10011110010010: Data_out <= 16'hA964	;
				14'b10011110010011: Data_out <= 16'hA95B	;
				14'b10011110010100: Data_out <= 16'hA952	;
				14'b10011110010101: Data_out <= 16'hA948	;
				14'b10011110010110: Data_out <= 16'hA93F	;
				14'b10011110010111: Data_out <= 16'hA936	;
				14'b10011110011000: Data_out <= 16'hA92D	;
				14'b10011110011001: Data_out <= 16'hA923	;
				14'b10011110011010: Data_out <= 16'hA91A	;
				14'b10011110011011: Data_out <= 16'hA911	;
				14'b10011110011100: Data_out <= 16'hA908	;
				14'b10011110011101: Data_out <= 16'hA8FE	;
				14'b10011110011110: Data_out <= 16'hA8F5	;
				14'b10011110011111: Data_out <= 16'hA8EC	;
				14'b10011110100000: Data_out <= 16'hA8E3	;
				14'b10011110100001: Data_out <= 16'hA8DA	;
				14'b10011110100010: Data_out <= 16'hA8D0	;
				14'b10011110100011: Data_out <= 16'hA8C7	;
				14'b10011110100100: Data_out <= 16'hA8BE	;
				14'b10011110100101: Data_out <= 16'hA8B5	;
				14'b10011110100110: Data_out <= 16'hA8AC	;
				14'b10011110100111: Data_out <= 16'hA8A2	;
				14'b10011110101000: Data_out <= 16'hA899	;
				14'b10011110101001: Data_out <= 16'hA890	;
				14'b10011110101010: Data_out <= 16'hA887	;
				14'b10011110101011: Data_out <= 16'hA87E	;
				14'b10011110101100: Data_out <= 16'hA875	;
				14'b10011110101101: Data_out <= 16'hA86B	;
				14'b10011110101110: Data_out <= 16'hA862	;
				14'b10011110101111: Data_out <= 16'hA859	;
				14'b10011110110000: Data_out <= 16'hA850	;
				14'b10011110110001: Data_out <= 16'hA847	;
				14'b10011110110010: Data_out <= 16'hA83E	;
				14'b10011110110011: Data_out <= 16'hA835	;
				14'b10011110110100: Data_out <= 16'hA82B	;
				14'b10011110110101: Data_out <= 16'hA822	;
				14'b10011110110110: Data_out <= 16'hA819	;
				14'b10011110110111: Data_out <= 16'hA810	;
				14'b10011110111000: Data_out <= 16'hA807	;
				14'b10011110111001: Data_out <= 16'hA7FE	;
				14'b10011110111010: Data_out <= 16'hA7F5	;
				14'b10011110111011: Data_out <= 16'hA7EB	;
				14'b10011110111100: Data_out <= 16'hA7E2	;
				14'b10011110111101: Data_out <= 16'hA7D9	;
				14'b10011110111110: Data_out <= 16'hA7D0	;
				14'b10011110111111: Data_out <= 16'hA7C7	;
				14'b10011111000000: Data_out <= 16'hA7BE	;
				14'b10011111000001: Data_out <= 16'hA7B5	;
				14'b10011111000010: Data_out <= 16'hA7AC	;
				14'b10011111000011: Data_out <= 16'hA7A3	;
				14'b10011111000100: Data_out <= 16'hA79A	;
				14'b10011111000101: Data_out <= 16'hA790	;
				14'b10011111000110: Data_out <= 16'hA787	;
				14'b10011111000111: Data_out <= 16'hA77E	;
				14'b10011111001000: Data_out <= 16'hA775	;
				14'b10011111001001: Data_out <= 16'hA76C	;
				14'b10011111001010: Data_out <= 16'hA763	;
				14'b10011111001011: Data_out <= 16'hA75A	;
				14'b10011111001100: Data_out <= 16'hA751	;
				14'b10011111001101: Data_out <= 16'hA748	;
				14'b10011111001110: Data_out <= 16'hA73F	;
				14'b10011111001111: Data_out <= 16'hA736	;
				14'b10011111010000: Data_out <= 16'hA72D	;
				14'b10011111010001: Data_out <= 16'hA724	;
				14'b10011111010010: Data_out <= 16'hA71B	;
				14'b10011111010011: Data_out <= 16'hA712	;
				14'b10011111010100: Data_out <= 16'hA709	;
				14'b10011111010101: Data_out <= 16'hA700	;
				14'b10011111010110: Data_out <= 16'hA6F7	;
				14'b10011111010111: Data_out <= 16'hA6ED	;
				14'b10011111011000: Data_out <= 16'hA6E4	;
				14'b10011111011001: Data_out <= 16'hA6DB	;
				14'b10011111011010: Data_out <= 16'hA6D2	;
				14'b10011111011011: Data_out <= 16'hA6C9	;
				14'b10011111011100: Data_out <= 16'hA6C0	;
				14'b10011111011101: Data_out <= 16'hA6B7	;
				14'b10011111011110: Data_out <= 16'hA6AE	;
				14'b10011111011111: Data_out <= 16'hA6A5	;
				14'b10011111100000: Data_out <= 16'hA69C	;
				14'b10011111100001: Data_out <= 16'hA693	;
				14'b10011111100010: Data_out <= 16'hA68A	;
				14'b10011111100011: Data_out <= 16'hA681	;
				14'b10011111100100: Data_out <= 16'hA678	;
				14'b10011111100101: Data_out <= 16'hA66F	;
				14'b10011111100110: Data_out <= 16'hA667	;
				14'b10011111100111: Data_out <= 16'hA65E	;
				14'b10011111101000: Data_out <= 16'hA655	;
				14'b10011111101001: Data_out <= 16'hA64C	;
				14'b10011111101010: Data_out <= 16'hA643	;
				14'b10011111101011: Data_out <= 16'hA63A	;
				14'b10011111101100: Data_out <= 16'hA631	;
				14'b10011111101101: Data_out <= 16'hA628	;
				14'b10011111101110: Data_out <= 16'hA61F	;
				14'b10011111101111: Data_out <= 16'hA616	;
				14'b10011111110000: Data_out <= 16'hA60D	;
				14'b10011111110001: Data_out <= 16'hA604	;
				14'b10011111110010: Data_out <= 16'hA5FB	;
				14'b10011111110011: Data_out <= 16'hA5F2	;
				14'b10011111110100: Data_out <= 16'hA5E9	;
				14'b10011111110101: Data_out <= 16'hA5E0	;
				14'b10011111110110: Data_out <= 16'hA5D7	;
				14'b10011111110111: Data_out <= 16'hA5CE	;
				14'b10011111111000: Data_out <= 16'hA5C6	;
				14'b10011111111001: Data_out <= 16'hA5BD	;
				14'b10011111111010: Data_out <= 16'hA5B4	;
				14'b10011111111011: Data_out <= 16'hA5AB	;
				14'b10011111111100: Data_out <= 16'hA5A2	;
				14'b10011111111101: Data_out <= 16'hA599	;
				14'b10011111111110: Data_out <= 16'hA590	;
				14'b10011111111111: Data_out <= 16'hA587	;
				14'b10100000000000: Data_out <= 16'hA57E	;
				14'b10100000000001: Data_out <= 16'hA575	;
				14'b10100000000010: Data_out <= 16'hA56D	;
				14'b10100000000011: Data_out <= 16'hA564	;
				14'b10100000000100: Data_out <= 16'hA55B	;
				14'b10100000000101: Data_out <= 16'hA552	;
				14'b10100000000110: Data_out <= 16'hA549	;
				14'b10100000000111: Data_out <= 16'hA540	;
				14'b10100000001000: Data_out <= 16'hA537	;
				14'b10100000001001: Data_out <= 16'hA52F	;
				14'b10100000001010: Data_out <= 16'hA526	;
				14'b10100000001011: Data_out <= 16'hA51D	;
				14'b10100000001100: Data_out <= 16'hA514	;
				14'b10100000001101: Data_out <= 16'hA50B	;
				14'b10100000001110: Data_out <= 16'hA502	;
				14'b10100000001111: Data_out <= 16'hA4F9	;
				14'b10100000010000: Data_out <= 16'hA4F1	;
				14'b10100000010001: Data_out <= 16'hA4E8	;
				14'b10100000010010: Data_out <= 16'hA4DF	;
				14'b10100000010011: Data_out <= 16'hA4D6	;
				14'b10100000010100: Data_out <= 16'hA4CD	;
				14'b10100000010101: Data_out <= 16'hA4C4	;
				14'b10100000010110: Data_out <= 16'hA4BC	;
				14'b10100000010111: Data_out <= 16'hA4B3	;
				14'b10100000011000: Data_out <= 16'hA4AA	;
				14'b10100000011001: Data_out <= 16'hA4A1	;
				14'b10100000011010: Data_out <= 16'hA498	;
				14'b10100000011011: Data_out <= 16'hA490	;
				14'b10100000011100: Data_out <= 16'hA487	;
				14'b10100000011101: Data_out <= 16'hA47E	;
				14'b10100000011110: Data_out <= 16'hA475	;
				14'b10100000011111: Data_out <= 16'hA46D	;
				14'b10100000100000: Data_out <= 16'hA464	;
				14'b10100000100001: Data_out <= 16'hA45B	;
				14'b10100000100010: Data_out <= 16'hA452	;
				14'b10100000100011: Data_out <= 16'hA449	;
				14'b10100000100100: Data_out <= 16'hA441	;
				14'b10100000100101: Data_out <= 16'hA438	;
				14'b10100000100110: Data_out <= 16'hA42F	;
				14'b10100000100111: Data_out <= 16'hA426	;
				14'b10100000101000: Data_out <= 16'hA41E	;
				14'b10100000101001: Data_out <= 16'hA415	;
				14'b10100000101010: Data_out <= 16'hA40C	;
				14'b10100000101011: Data_out <= 16'hA403	;
				14'b10100000101100: Data_out <= 16'hA3FB	;
				14'b10100000101101: Data_out <= 16'hA3F2	;
				14'b10100000101110: Data_out <= 16'hA3E9	;
				14'b10100000101111: Data_out <= 16'hA3E0	;
				14'b10100000110000: Data_out <= 16'hA3D8	;
				14'b10100000110001: Data_out <= 16'hA3CF	;
				14'b10100000110010: Data_out <= 16'hA3C6	;
				14'b10100000110011: Data_out <= 16'hA3BE	;
				14'b10100000110100: Data_out <= 16'hA3B5	;
				14'b10100000110101: Data_out <= 16'hA3AC	;
				14'b10100000110110: Data_out <= 16'hA3A4	;
				14'b10100000110111: Data_out <= 16'hA39B	;
				14'b10100000111000: Data_out <= 16'hA392	;
				14'b10100000111001: Data_out <= 16'hA389	;
				14'b10100000111010: Data_out <= 16'hA381	;
				14'b10100000111011: Data_out <= 16'hA378	;
				14'b10100000111100: Data_out <= 16'hA36F	;
				14'b10100000111101: Data_out <= 16'hA367	;
				14'b10100000111110: Data_out <= 16'hA35E	;
				14'b10100000111111: Data_out <= 16'hA355	;
				14'b10100001000000: Data_out <= 16'hA34D	;
				14'b10100001000001: Data_out <= 16'hA344	;
				14'b10100001000010: Data_out <= 16'hA33B	;
				14'b10100001000011: Data_out <= 16'hA333	;
				14'b10100001000100: Data_out <= 16'hA32A	;
				14'b10100001000101: Data_out <= 16'hA321	;
				14'b10100001000110: Data_out <= 16'hA319	;
				14'b10100001000111: Data_out <= 16'hA310	;
				14'b10100001001000: Data_out <= 16'hA307	;
				14'b10100001001001: Data_out <= 16'hA2FF	;
				14'b10100001001010: Data_out <= 16'hA2F6	;
				14'b10100001001011: Data_out <= 16'hA2EE	;
				14'b10100001001100: Data_out <= 16'hA2E5	;
				14'b10100001001101: Data_out <= 16'hA2DC	;
				14'b10100001001110: Data_out <= 16'hA2D4	;
				14'b10100001001111: Data_out <= 16'hA2CB	;
				14'b10100001010000: Data_out <= 16'hA2C3	;
				14'b10100001010001: Data_out <= 16'hA2BA	;
				14'b10100001010010: Data_out <= 16'hA2B1	;
				14'b10100001010011: Data_out <= 16'hA2A9	;
				14'b10100001010100: Data_out <= 16'hA2A0	;
				14'b10100001010101: Data_out <= 16'hA298	;
				14'b10100001010110: Data_out <= 16'hA28F	;
				14'b10100001010111: Data_out <= 16'hA286	;
				14'b10100001011000: Data_out <= 16'hA27E	;
				14'b10100001011001: Data_out <= 16'hA275	;
				14'b10100001011010: Data_out <= 16'hA26D	;
				14'b10100001011011: Data_out <= 16'hA264	;
				14'b10100001011100: Data_out <= 16'hA25B	;
				14'b10100001011101: Data_out <= 16'hA253	;
				14'b10100001011110: Data_out <= 16'hA24A	;
				14'b10100001011111: Data_out <= 16'hA242	;
				14'b10100001100000: Data_out <= 16'hA239	;
				14'b10100001100001: Data_out <= 16'hA231	;
				14'b10100001100010: Data_out <= 16'hA228	;
				14'b10100001100011: Data_out <= 16'hA220	;
				14'b10100001100100: Data_out <= 16'hA217	;
				14'b10100001100101: Data_out <= 16'hA20E	;
				14'b10100001100110: Data_out <= 16'hA206	;
				14'b10100001100111: Data_out <= 16'hA1FD	;
				14'b10100001101000: Data_out <= 16'hA1F5	;
				14'b10100001101001: Data_out <= 16'hA1EC	;
				14'b10100001101010: Data_out <= 16'hA1E4	;
				14'b10100001101011: Data_out <= 16'hA1DB	;
				14'b10100001101100: Data_out <= 16'hA1D3	;
				14'b10100001101101: Data_out <= 16'hA1CA	;
				14'b10100001101110: Data_out <= 16'hA1C2	;
				14'b10100001101111: Data_out <= 16'hA1B9	;
				14'b10100001110000: Data_out <= 16'hA1B1	;
				14'b10100001110001: Data_out <= 16'hA1A8	;
				14'b10100001110010: Data_out <= 16'hA1A0	;
				14'b10100001110011: Data_out <= 16'hA197	;
				14'b10100001110100: Data_out <= 16'hA18F	;
				14'b10100001110101: Data_out <= 16'hA186	;
				14'b10100001110110: Data_out <= 16'hA17E	;
				14'b10100001110111: Data_out <= 16'hA175	;
				14'b10100001111000: Data_out <= 16'hA16D	;
				14'b10100001111001: Data_out <= 16'hA165	;
				14'b10100001111010: Data_out <= 16'hA15C	;
				14'b10100001111011: Data_out <= 16'hA154	;
				14'b10100001111100: Data_out <= 16'hA14B	;
				14'b10100001111101: Data_out <= 16'hA143	;
				14'b10100001111110: Data_out <= 16'hA13A	;
				14'b10100001111111: Data_out <= 16'hA132	;
				14'b10100010000000: Data_out <= 16'hA129	;
				14'b10100010000001: Data_out <= 16'hA121	;
				14'b10100010000010: Data_out <= 16'hA118	;
				14'b10100010000011: Data_out <= 16'hA110	;
				14'b10100010000100: Data_out <= 16'hA108	;
				14'b10100010000101: Data_out <= 16'hA0FF	;
				14'b10100010000110: Data_out <= 16'hA0F7	;
				14'b10100010000111: Data_out <= 16'hA0EE	;
				14'b10100010001000: Data_out <= 16'hA0E6	;
				14'b10100010001001: Data_out <= 16'hA0DE	;
				14'b10100010001010: Data_out <= 16'hA0D5	;
				14'b10100010001011: Data_out <= 16'hA0CD	;
				14'b10100010001100: Data_out <= 16'hA0C4	;
				14'b10100010001101: Data_out <= 16'hA0BC	;
				14'b10100010001110: Data_out <= 16'hA0B4	;
				14'b10100010001111: Data_out <= 16'hA0AB	;
				14'b10100010010000: Data_out <= 16'hA0A3	;
				14'b10100010010001: Data_out <= 16'hA09A	;
				14'b10100010010010: Data_out <= 16'hA092	;
				14'b10100010010011: Data_out <= 16'hA08A	;
				14'b10100010010100: Data_out <= 16'hA081	;
				14'b10100010010101: Data_out <= 16'hA079	;
				14'b10100010010110: Data_out <= 16'hA071	;
				14'b10100010010111: Data_out <= 16'hA068	;
				14'b10100010011000: Data_out <= 16'hA060	;
				14'b10100010011001: Data_out <= 16'hA058	;
				14'b10100010011010: Data_out <= 16'hA04F	;
				14'b10100010011011: Data_out <= 16'hA047	;
				14'b10100010011100: Data_out <= 16'hA03E	;
				14'b10100010011101: Data_out <= 16'hA036	;
				14'b10100010011110: Data_out <= 16'hA02E	;
				14'b10100010011111: Data_out <= 16'hA025	;
				14'b10100010100000: Data_out <= 16'hA01D	;
				14'b10100010100001: Data_out <= 16'hA015	;
				14'b10100010100010: Data_out <= 16'hA00D	;
				14'b10100010100011: Data_out <= 16'hA004	;
				14'b10100010100100: Data_out <= 16'h9FFC	;
				14'b10100010100101: Data_out <= 16'h9FF4	;
				14'b10100010100110: Data_out <= 16'h9FEB	;
				14'b10100010100111: Data_out <= 16'h9FE3	;
				14'b10100010101000: Data_out <= 16'h9FDB	;
				14'b10100010101001: Data_out <= 16'h9FD2	;
				14'b10100010101010: Data_out <= 16'h9FCA	;
				14'b10100010101011: Data_out <= 16'h9FC2	;
				14'b10100010101100: Data_out <= 16'h9FBA	;
				14'b10100010101101: Data_out <= 16'h9FB1	;
				14'b10100010101110: Data_out <= 16'h9FA9	;
				14'b10100010101111: Data_out <= 16'h9FA1	;
				14'b10100010110000: Data_out <= 16'h9F98	;
				14'b10100010110001: Data_out <= 16'h9F90	;
				14'b10100010110010: Data_out <= 16'h9F88	;
				14'b10100010110011: Data_out <= 16'h9F80	;
				14'b10100010110100: Data_out <= 16'h9F77	;
				14'b10100010110101: Data_out <= 16'h9F6F	;
				14'b10100010110110: Data_out <= 16'h9F67	;
				14'b10100010110111: Data_out <= 16'h9F5F	;
				14'b10100010111000: Data_out <= 16'h9F56	;
				14'b10100010111001: Data_out <= 16'h9F4E	;
				14'b10100010111010: Data_out <= 16'h9F46	;
				14'b10100010111011: Data_out <= 16'h9F3E	;
				14'b10100010111100: Data_out <= 16'h9F35	;
				14'b10100010111101: Data_out <= 16'h9F2D	;
				14'b10100010111110: Data_out <= 16'h9F25	;
				14'b10100010111111: Data_out <= 16'h9F1D	;
				14'b10100011000000: Data_out <= 16'h9F15	;
				14'b10100011000001: Data_out <= 16'h9F0C	;
				14'b10100011000010: Data_out <= 16'h9F04	;
				14'b10100011000011: Data_out <= 16'h9EFC	;
				14'b10100011000100: Data_out <= 16'h9EF4	;
				14'b10100011000101: Data_out <= 16'h9EEC	;
				14'b10100011000110: Data_out <= 16'h9EE3	;
				14'b10100011000111: Data_out <= 16'h9EDB	;
				14'b10100011001000: Data_out <= 16'h9ED3	;
				14'b10100011001001: Data_out <= 16'h9ECB	;
				14'b10100011001010: Data_out <= 16'h9EC3	;
				14'b10100011001011: Data_out <= 16'h9EBB	;
				14'b10100011001100: Data_out <= 16'h9EB2	;
				14'b10100011001101: Data_out <= 16'h9EAA	;
				14'b10100011001110: Data_out <= 16'h9EA2	;
				14'b10100011001111: Data_out <= 16'h9E9A	;
				14'b10100011010000: Data_out <= 16'h9E92	;
				14'b10100011010001: Data_out <= 16'h9E8A	;
				14'b10100011010010: Data_out <= 16'h9E81	;
				14'b10100011010011: Data_out <= 16'h9E79	;
				14'b10100011010100: Data_out <= 16'h9E71	;
				14'b10100011010101: Data_out <= 16'h9E69	;
				14'b10100011010110: Data_out <= 16'h9E61	;
				14'b10100011010111: Data_out <= 16'h9E59	;
				14'b10100011011000: Data_out <= 16'h9E51	;
				14'b10100011011001: Data_out <= 16'h9E49	;
				14'b10100011011010: Data_out <= 16'h9E40	;
				14'b10100011011011: Data_out <= 16'h9E38	;
				14'b10100011011100: Data_out <= 16'h9E30	;
				14'b10100011011101: Data_out <= 16'h9E28	;
				14'b10100011011110: Data_out <= 16'h9E20	;
				14'b10100011011111: Data_out <= 16'h9E18	;
				14'b10100011100000: Data_out <= 16'h9E10	;
				14'b10100011100001: Data_out <= 16'h9E08	;
				14'b10100011100010: Data_out <= 16'h9E00	;
				14'b10100011100011: Data_out <= 16'h9DF8	;
				14'b10100011100100: Data_out <= 16'h9DF0	;
				14'b10100011100101: Data_out <= 16'h9DE7	;
				14'b10100011100110: Data_out <= 16'h9DDF	;
				14'b10100011100111: Data_out <= 16'h9DD7	;
				14'b10100011101000: Data_out <= 16'h9DCF	;
				14'b10100011101001: Data_out <= 16'h9DC7	;
				14'b10100011101010: Data_out <= 16'h9DBF	;
				14'b10100011101011: Data_out <= 16'h9DB7	;
				14'b10100011101100: Data_out <= 16'h9DAF	;
				14'b10100011101101: Data_out <= 16'h9DA7	;
				14'b10100011101110: Data_out <= 16'h9D9F	;
				14'b10100011101111: Data_out <= 16'h9D97	;
				14'b10100011110000: Data_out <= 16'h9D8F	;
				14'b10100011110001: Data_out <= 16'h9D87	;
				14'b10100011110010: Data_out <= 16'h9D7F	;
				14'b10100011110011: Data_out <= 16'h9D77	;
				14'b10100011110100: Data_out <= 16'h9D6F	;
				14'b10100011110101: Data_out <= 16'h9D67	;
				14'b10100011110110: Data_out <= 16'h9D5F	;
				14'b10100011110111: Data_out <= 16'h9D57	;
				14'b10100011111000: Data_out <= 16'h9D4F	;
				14'b10100011111001: Data_out <= 16'h9D47	;
				14'b10100011111010: Data_out <= 16'h9D3F	;
				14'b10100011111011: Data_out <= 16'h9D37	;
				14'b10100011111100: Data_out <= 16'h9D2F	;
				14'b10100011111101: Data_out <= 16'h9D27	;
				14'b10100011111110: Data_out <= 16'h9D1F	;
				14'b10100011111111: Data_out <= 16'h9D17	;
				14'b10100100000000: Data_out <= 16'h9D0F	;
				14'b10100100000001: Data_out <= 16'h9D07	;
				14'b10100100000010: Data_out <= 16'h9CFF	;
				14'b10100100000011: Data_out <= 16'h9CF7	;
				14'b10100100000100: Data_out <= 16'h9CEF	;
				14'b10100100000101: Data_out <= 16'h9CE7	;
				14'b10100100000110: Data_out <= 16'h9CDF	;
				14'b10100100000111: Data_out <= 16'h9CD7	;
				14'b10100100001000: Data_out <= 16'h9CCF	;
				14'b10100100001001: Data_out <= 16'h9CC7	;
				14'b10100100001010: Data_out <= 16'h9CBF	;
				14'b10100100001011: Data_out <= 16'h9CB7	;
				14'b10100100001100: Data_out <= 16'h9CAF	;
				14'b10100100001101: Data_out <= 16'h9CA8	;
				14'b10100100001110: Data_out <= 16'h9CA0	;
				14'b10100100001111: Data_out <= 16'h9C98	;
				14'b10100100010000: Data_out <= 16'h9C90	;
				14'b10100100010001: Data_out <= 16'h9C88	;
				14'b10100100010010: Data_out <= 16'h9C80	;
				14'b10100100010011: Data_out <= 16'h9C78	;
				14'b10100100010100: Data_out <= 16'h9C70	;
				14'b10100100010101: Data_out <= 16'h9C68	;
				14'b10100100010110: Data_out <= 16'h9C60	;
				14'b10100100010111: Data_out <= 16'h9C59	;
				14'b10100100011000: Data_out <= 16'h9C51	;
				14'b10100100011001: Data_out <= 16'h9C49	;
				14'b10100100011010: Data_out <= 16'h9C41	;
				14'b10100100011011: Data_out <= 16'h9C39	;
				14'b10100100011100: Data_out <= 16'h9C31	;
				14'b10100100011101: Data_out <= 16'h9C29	;
				14'b10100100011110: Data_out <= 16'h9C21	;
				14'b10100100011111: Data_out <= 16'h9C1A	;
				14'b10100100100000: Data_out <= 16'h9C12	;
				14'b10100100100001: Data_out <= 16'h9C0A	;
				14'b10100100100010: Data_out <= 16'h9C02	;
				14'b10100100100011: Data_out <= 16'h9BFA	;
				14'b10100100100100: Data_out <= 16'h9BF2	;
				14'b10100100100101: Data_out <= 16'h9BEA	;
				14'b10100100100110: Data_out <= 16'h9BE3	;
				14'b10100100100111: Data_out <= 16'h9BDB	;
				14'b10100100101000: Data_out <= 16'h9BD3	;
				14'b10100100101001: Data_out <= 16'h9BCB	;
				14'b10100100101010: Data_out <= 16'h9BC3	;
				14'b10100100101011: Data_out <= 16'h9BBC	;
				14'b10100100101100: Data_out <= 16'h9BB4	;
				14'b10100100101101: Data_out <= 16'h9BAC	;
				14'b10100100101110: Data_out <= 16'h9BA4	;
				14'b10100100101111: Data_out <= 16'h9B9C	;
				14'b10100100110000: Data_out <= 16'h9B95	;
				14'b10100100110001: Data_out <= 16'h9B8D	;
				14'b10100100110010: Data_out <= 16'h9B85	;
				14'b10100100110011: Data_out <= 16'h9B7D	;
				14'b10100100110100: Data_out <= 16'h9B75	;
				14'b10100100110101: Data_out <= 16'h9B6E	;
				14'b10100100110110: Data_out <= 16'h9B66	;
				14'b10100100110111: Data_out <= 16'h9B5E	;
				14'b10100100111000: Data_out <= 16'h9B56	;
				14'b10100100111001: Data_out <= 16'h9B4F	;
				14'b10100100111010: Data_out <= 16'h9B47	;
				14'b10100100111011: Data_out <= 16'h9B3F	;
				14'b10100100111100: Data_out <= 16'h9B37	;
				14'b10100100111101: Data_out <= 16'h9B30	;
				14'b10100100111110: Data_out <= 16'h9B28	;
				14'b10100100111111: Data_out <= 16'h9B20	;
				14'b10100101000000: Data_out <= 16'h9B18	;
				14'b10100101000001: Data_out <= 16'h9B11	;
				14'b10100101000010: Data_out <= 16'h9B09	;
				14'b10100101000011: Data_out <= 16'h9B01	;
				14'b10100101000100: Data_out <= 16'h9AF9	;
				14'b10100101000101: Data_out <= 16'h9AF2	;
				14'b10100101000110: Data_out <= 16'h9AEA	;
				14'b10100101000111: Data_out <= 16'h9AE2	;
				14'b10100101001000: Data_out <= 16'h9ADB	;
				14'b10100101001001: Data_out <= 16'h9AD3	;
				14'b10100101001010: Data_out <= 16'h9ACB	;
				14'b10100101001011: Data_out <= 16'h9AC4	;
				14'b10100101001100: Data_out <= 16'h9ABC	;
				14'b10100101001101: Data_out <= 16'h9AB4	;
				14'b10100101001110: Data_out <= 16'h9AAC	;
				14'b10100101001111: Data_out <= 16'h9AA5	;
				14'b10100101010000: Data_out <= 16'h9A9D	;
				14'b10100101010001: Data_out <= 16'h9A95	;
				14'b10100101010010: Data_out <= 16'h9A8E	;
				14'b10100101010011: Data_out <= 16'h9A86	;
				14'b10100101010100: Data_out <= 16'h9A7E	;
				14'b10100101010101: Data_out <= 16'h9A77	;
				14'b10100101010110: Data_out <= 16'h9A6F	;
				14'b10100101010111: Data_out <= 16'h9A68	;
				14'b10100101011000: Data_out <= 16'h9A60	;
				14'b10100101011001: Data_out <= 16'h9A58	;
				14'b10100101011010: Data_out <= 16'h9A51	;
				14'b10100101011011: Data_out <= 16'h9A49	;
				14'b10100101011100: Data_out <= 16'h9A41	;
				14'b10100101011101: Data_out <= 16'h9A3A	;
				14'b10100101011110: Data_out <= 16'h9A32	;
				14'b10100101011111: Data_out <= 16'h9A2B	;
				14'b10100101100000: Data_out <= 16'h9A23	;
				14'b10100101100001: Data_out <= 16'h9A1B	;
				14'b10100101100010: Data_out <= 16'h9A14	;
				14'b10100101100011: Data_out <= 16'h9A0C	;
				14'b10100101100100: Data_out <= 16'h9A05	;
				14'b10100101100101: Data_out <= 16'h99FD	;
				14'b10100101100110: Data_out <= 16'h99F5	;
				14'b10100101100111: Data_out <= 16'h99EE	;
				14'b10100101101000: Data_out <= 16'h99E6	;
				14'b10100101101001: Data_out <= 16'h99DF	;
				14'b10100101101010: Data_out <= 16'h99D7	;
				14'b10100101101011: Data_out <= 16'h99CF	;
				14'b10100101101100: Data_out <= 16'h99C8	;
				14'b10100101101101: Data_out <= 16'h99C0	;
				14'b10100101101110: Data_out <= 16'h99B9	;
				14'b10100101101111: Data_out <= 16'h99B1	;
				14'b10100101110000: Data_out <= 16'h99AA	;
				14'b10100101110001: Data_out <= 16'h99A2	;
				14'b10100101110010: Data_out <= 16'h999B	;
				14'b10100101110011: Data_out <= 16'h9993	;
				14'b10100101110100: Data_out <= 16'h998C	;
				14'b10100101110101: Data_out <= 16'h9984	;
				14'b10100101110110: Data_out <= 16'h997C	;
				14'b10100101110111: Data_out <= 16'h9975	;
				14'b10100101111000: Data_out <= 16'h996D	;
				14'b10100101111001: Data_out <= 16'h9966	;
				14'b10100101111010: Data_out <= 16'h995E	;
				14'b10100101111011: Data_out <= 16'h9957	;
				14'b10100101111100: Data_out <= 16'h994F	;
				14'b10100101111101: Data_out <= 16'h9948	;
				14'b10100101111110: Data_out <= 16'h9940	;
				14'b10100101111111: Data_out <= 16'h9939	;
				14'b10100110000000: Data_out <= 16'h9931	;
				14'b10100110000001: Data_out <= 16'h992A	;
				14'b10100110000010: Data_out <= 16'h9922	;
				14'b10100110000011: Data_out <= 16'h991B	;
				14'b10100110000100: Data_out <= 16'h9913	;
				14'b10100110000101: Data_out <= 16'h990C	;
				14'b10100110000110: Data_out <= 16'h9905	;
				14'b10100110000111: Data_out <= 16'h98FD	;
				14'b10100110001000: Data_out <= 16'h98F6	;
				14'b10100110001001: Data_out <= 16'h98EE	;
				14'b10100110001010: Data_out <= 16'h98E7	;
				14'b10100110001011: Data_out <= 16'h98DF	;
				14'b10100110001100: Data_out <= 16'h98D8	;
				14'b10100110001101: Data_out <= 16'h98D0	;
				14'b10100110001110: Data_out <= 16'h98C9	;
				14'b10100110001111: Data_out <= 16'h98C2	;
				14'b10100110010000: Data_out <= 16'h98BA	;
				14'b10100110010001: Data_out <= 16'h98B3	;
				14'b10100110010010: Data_out <= 16'h98AB	;
				14'b10100110010011: Data_out <= 16'h98A4	;
				14'b10100110010100: Data_out <= 16'h989C	;
				14'b10100110010101: Data_out <= 16'h9895	;
				14'b10100110010110: Data_out <= 16'h988E	;
				14'b10100110010111: Data_out <= 16'h9886	;
				14'b10100110011000: Data_out <= 16'h987F	;
				14'b10100110011001: Data_out <= 16'h9877	;
				14'b10100110011010: Data_out <= 16'h9870	;
				14'b10100110011011: Data_out <= 16'h9869	;
				14'b10100110011100: Data_out <= 16'h9861	;
				14'b10100110011101: Data_out <= 16'h985A	;
				14'b10100110011110: Data_out <= 16'h9853	;
				14'b10100110011111: Data_out <= 16'h984B	;
				14'b10100110100000: Data_out <= 16'h9844	;
				14'b10100110100001: Data_out <= 16'h983C	;
				14'b10100110100010: Data_out <= 16'h9835	;
				14'b10100110100011: Data_out <= 16'h982E	;
				14'b10100110100100: Data_out <= 16'h9826	;
				14'b10100110100101: Data_out <= 16'h981F	;
				14'b10100110100110: Data_out <= 16'h9818	;
				14'b10100110100111: Data_out <= 16'h9810	;
				14'b10100110101000: Data_out <= 16'h9809	;
				14'b10100110101001: Data_out <= 16'h9802	;
				14'b10100110101010: Data_out <= 16'h97FA	;
				14'b10100110101011: Data_out <= 16'h97F3	;
				14'b10100110101100: Data_out <= 16'h97EC	;
				14'b10100110101101: Data_out <= 16'h97E4	;
				14'b10100110101110: Data_out <= 16'h97DD	;
				14'b10100110101111: Data_out <= 16'h97D6	;
				14'b10100110110000: Data_out <= 16'h97CF	;
				14'b10100110110001: Data_out <= 16'h97C7	;
				14'b10100110110010: Data_out <= 16'h97C0	;
				14'b10100110110011: Data_out <= 16'h97B9	;
				14'b10100110110100: Data_out <= 16'h97B1	;
				14'b10100110110101: Data_out <= 16'h97AA	;
				14'b10100110110110: Data_out <= 16'h97A3	;
				14'b10100110110111: Data_out <= 16'h979C	;
				14'b10100110111000: Data_out <= 16'h9794	;
				14'b10100110111001: Data_out <= 16'h978D	;
				14'b10100110111010: Data_out <= 16'h9786	;
				14'b10100110111011: Data_out <= 16'h977F	;
				14'b10100110111100: Data_out <= 16'h9777	;
				14'b10100110111101: Data_out <= 16'h9770	;
				14'b10100110111110: Data_out <= 16'h9769	;
				14'b10100110111111: Data_out <= 16'h9762	;
				14'b10100111000000: Data_out <= 16'h975A	;
				14'b10100111000001: Data_out <= 16'h9753	;
				14'b10100111000010: Data_out <= 16'h974C	;
				14'b10100111000011: Data_out <= 16'h9745	;
				14'b10100111000100: Data_out <= 16'h973D	;
				14'b10100111000101: Data_out <= 16'h9736	;
				14'b10100111000110: Data_out <= 16'h972F	;
				14'b10100111000111: Data_out <= 16'h9728	;
				14'b10100111001000: Data_out <= 16'h9721	;
				14'b10100111001001: Data_out <= 16'h9719	;
				14'b10100111001010: Data_out <= 16'h9712	;
				14'b10100111001011: Data_out <= 16'h970B	;
				14'b10100111001100: Data_out <= 16'h9704	;
				14'b10100111001101: Data_out <= 16'h96FD	;
				14'b10100111001110: Data_out <= 16'h96F5	;
				14'b10100111001111: Data_out <= 16'h96EE	;
				14'b10100111010000: Data_out <= 16'h96E7	;
				14'b10100111010001: Data_out <= 16'h96E0	;
				14'b10100111010010: Data_out <= 16'h96D9	;
				14'b10100111010011: Data_out <= 16'h96D2	;
				14'b10100111010100: Data_out <= 16'h96CA	;
				14'b10100111010101: Data_out <= 16'h96C3	;
				14'b10100111010110: Data_out <= 16'h96BC	;
				14'b10100111010111: Data_out <= 16'h96B5	;
				14'b10100111011000: Data_out <= 16'h96AE	;
				14'b10100111011001: Data_out <= 16'h96A7	;
				14'b10100111011010: Data_out <= 16'h96A0	;
				14'b10100111011011: Data_out <= 16'h9698	;
				14'b10100111011100: Data_out <= 16'h9691	;
				14'b10100111011101: Data_out <= 16'h968A	;
				14'b10100111011110: Data_out <= 16'h9683	;
				14'b10100111011111: Data_out <= 16'h967C	;
				14'b10100111100000: Data_out <= 16'h9675	;
				14'b10100111100001: Data_out <= 16'h966E	;
				14'b10100111100010: Data_out <= 16'h9667	;
				14'b10100111100011: Data_out <= 16'h965F	;
				14'b10100111100100: Data_out <= 16'h9658	;
				14'b10100111100101: Data_out <= 16'h9651	;
				14'b10100111100110: Data_out <= 16'h964A	;
				14'b10100111100111: Data_out <= 16'h9643	;
				14'b10100111101000: Data_out <= 16'h963C	;
				14'b10100111101001: Data_out <= 16'h9635	;
				14'b10100111101010: Data_out <= 16'h962E	;
				14'b10100111101011: Data_out <= 16'h9627	;
				14'b10100111101100: Data_out <= 16'h9620	;
				14'b10100111101101: Data_out <= 16'h9619	;
				14'b10100111101110: Data_out <= 16'h9612	;
				14'b10100111101111: Data_out <= 16'h960B	;
				14'b10100111110000: Data_out <= 16'h9604	;
				14'b10100111110001: Data_out <= 16'h95FD	;
				14'b10100111110010: Data_out <= 16'h95F5	;
				14'b10100111110011: Data_out <= 16'h95EE	;
				14'b10100111110100: Data_out <= 16'h95E7	;
				14'b10100111110101: Data_out <= 16'h95E0	;
				14'b10100111110110: Data_out <= 16'h95D9	;
				14'b10100111110111: Data_out <= 16'h95D2	;
				14'b10100111111000: Data_out <= 16'h95CB	;
				14'b10100111111001: Data_out <= 16'h95C4	;
				14'b10100111111010: Data_out <= 16'h95BD	;
				14'b10100111111011: Data_out <= 16'h95B6	;
				14'b10100111111100: Data_out <= 16'h95AF	;
				14'b10100111111101: Data_out <= 16'h95A8	;
				14'b10100111111110: Data_out <= 16'h95A1	;
				14'b10100111111111: Data_out <= 16'h959A	;
				14'b10101000000000: Data_out <= 16'h9593	;
				14'b10101000000001: Data_out <= 16'h958C	;
				14'b10101000000010: Data_out <= 16'h9585	;
				14'b10101000000011: Data_out <= 16'h957E	;
				14'b10101000000100: Data_out <= 16'h9577	;
				14'b10101000000101: Data_out <= 16'h9570	;
				14'b10101000000110: Data_out <= 16'h956A	;
				14'b10101000000111: Data_out <= 16'h9563	;
				14'b10101000001000: Data_out <= 16'h955C	;
				14'b10101000001001: Data_out <= 16'h9555	;
				14'b10101000001010: Data_out <= 16'h954E	;
				14'b10101000001011: Data_out <= 16'h9547	;
				14'b10101000001100: Data_out <= 16'h9540	;
				14'b10101000001101: Data_out <= 16'h9539	;
				14'b10101000001110: Data_out <= 16'h9532	;
				14'b10101000001111: Data_out <= 16'h952B	;
				14'b10101000010000: Data_out <= 16'h9524	;
				14'b10101000010001: Data_out <= 16'h951D	;
				14'b10101000010010: Data_out <= 16'h9516	;
				14'b10101000010011: Data_out <= 16'h950F	;
				14'b10101000010100: Data_out <= 16'h9509	;
				14'b10101000010101: Data_out <= 16'h9502	;
				14'b10101000010110: Data_out <= 16'h94FB	;
				14'b10101000010111: Data_out <= 16'h94F4	;
				14'b10101000011000: Data_out <= 16'h94ED	;
				14'b10101000011001: Data_out <= 16'h94E6	;
				14'b10101000011010: Data_out <= 16'h94DF	;
				14'b10101000011011: Data_out <= 16'h94D8	;
				14'b10101000011100: Data_out <= 16'h94D1	;
				14'b10101000011101: Data_out <= 16'h94CB	;
				14'b10101000011110: Data_out <= 16'h94C4	;
				14'b10101000011111: Data_out <= 16'h94BD	;
				14'b10101000100000: Data_out <= 16'h94B6	;
				14'b10101000100001: Data_out <= 16'h94AF	;
				14'b10101000100010: Data_out <= 16'h94A8	;
				14'b10101000100011: Data_out <= 16'h94A1	;
				14'b10101000100100: Data_out <= 16'h949B	;
				14'b10101000100101: Data_out <= 16'h9494	;
				14'b10101000100110: Data_out <= 16'h948D	;
				14'b10101000100111: Data_out <= 16'h9486	;
				14'b10101000101000: Data_out <= 16'h947F	;
				14'b10101000101001: Data_out <= 16'h9478	;
				14'b10101000101010: Data_out <= 16'h9472	;
				14'b10101000101011: Data_out <= 16'h946B	;
				14'b10101000101100: Data_out <= 16'h9464	;
				14'b10101000101101: Data_out <= 16'h945D	;
				14'b10101000101110: Data_out <= 16'h9456	;
				14'b10101000101111: Data_out <= 16'h9450	;
				14'b10101000110000: Data_out <= 16'h9449	;
				14'b10101000110001: Data_out <= 16'h9442	;
				14'b10101000110010: Data_out <= 16'h943B	;
				14'b10101000110011: Data_out <= 16'h9435	;
				14'b10101000110100: Data_out <= 16'h942E	;
				14'b10101000110101: Data_out <= 16'h9427	;
				14'b10101000110110: Data_out <= 16'h9420	;
				14'b10101000110111: Data_out <= 16'h9419	;
				14'b10101000111000: Data_out <= 16'h9413	;
				14'b10101000111001: Data_out <= 16'h940C	;
				14'b10101000111010: Data_out <= 16'h9405	;
				14'b10101000111011: Data_out <= 16'h93FE	;
				14'b10101000111100: Data_out <= 16'h93F8	;
				14'b10101000111101: Data_out <= 16'h93F1	;
				14'b10101000111110: Data_out <= 16'h93EA	;
				14'b10101000111111: Data_out <= 16'h93E4	;
				14'b10101001000000: Data_out <= 16'h93DD	;
				14'b10101001000001: Data_out <= 16'h93D6	;
				14'b10101001000010: Data_out <= 16'h93CF	;
				14'b10101001000011: Data_out <= 16'h93C9	;
				14'b10101001000100: Data_out <= 16'h93C2	;
				14'b10101001000101: Data_out <= 16'h93BB	;
				14'b10101001000110: Data_out <= 16'h93B5	;
				14'b10101001000111: Data_out <= 16'h93AE	;
				14'b10101001001000: Data_out <= 16'h93A7	;
				14'b10101001001001: Data_out <= 16'h93A0	;
				14'b10101001001010: Data_out <= 16'h939A	;
				14'b10101001001011: Data_out <= 16'h9393	;
				14'b10101001001100: Data_out <= 16'h938C	;
				14'b10101001001101: Data_out <= 16'h9386	;
				14'b10101001001110: Data_out <= 16'h937F	;
				14'b10101001001111: Data_out <= 16'h9378	;
				14'b10101001010000: Data_out <= 16'h9372	;
				14'b10101001010001: Data_out <= 16'h936B	;
				14'b10101001010010: Data_out <= 16'h9364	;
				14'b10101001010011: Data_out <= 16'h935E	;
				14'b10101001010100: Data_out <= 16'h9357	;
				14'b10101001010101: Data_out <= 16'h9351	;
				14'b10101001010110: Data_out <= 16'h934A	;
				14'b10101001010111: Data_out <= 16'h9343	;
				14'b10101001011000: Data_out <= 16'h933D	;
				14'b10101001011001: Data_out <= 16'h9336	;
				14'b10101001011010: Data_out <= 16'h932F	;
				14'b10101001011011: Data_out <= 16'h9329	;
				14'b10101001011100: Data_out <= 16'h9322	;
				14'b10101001011101: Data_out <= 16'h931C	;
				14'b10101001011110: Data_out <= 16'h9315	;
				14'b10101001011111: Data_out <= 16'h930E	;
				14'b10101001100000: Data_out <= 16'h9308	;
				14'b10101001100001: Data_out <= 16'h9301	;
				14'b10101001100010: Data_out <= 16'h92FB	;
				14'b10101001100011: Data_out <= 16'h92F4	;
				14'b10101001100100: Data_out <= 16'h92ED	;
				14'b10101001100101: Data_out <= 16'h92E7	;
				14'b10101001100110: Data_out <= 16'h92E0	;
				14'b10101001100111: Data_out <= 16'h92DA	;
				14'b10101001101000: Data_out <= 16'h92D3	;
				14'b10101001101001: Data_out <= 16'h92CD	;
				14'b10101001101010: Data_out <= 16'h92C6	;
				14'b10101001101011: Data_out <= 16'h92BF	;
				14'b10101001101100: Data_out <= 16'h92B9	;
				14'b10101001101101: Data_out <= 16'h92B2	;
				14'b10101001101110: Data_out <= 16'h92AC	;
				14'b10101001101111: Data_out <= 16'h92A5	;
				14'b10101001110000: Data_out <= 16'h929F	;
				14'b10101001110001: Data_out <= 16'h9298	;
				14'b10101001110010: Data_out <= 16'h9292	;
				14'b10101001110011: Data_out <= 16'h928B	;
				14'b10101001110100: Data_out <= 16'h9285	;
				14'b10101001110101: Data_out <= 16'h927E	;
				14'b10101001110110: Data_out <= 16'h9278	;
				14'b10101001110111: Data_out <= 16'h9271	;
				14'b10101001111000: Data_out <= 16'h926B	;
				14'b10101001111001: Data_out <= 16'h9264	;
				14'b10101001111010: Data_out <= 16'h925E	;
				14'b10101001111011: Data_out <= 16'h9257	;
				14'b10101001111100: Data_out <= 16'h9251	;
				14'b10101001111101: Data_out <= 16'h924A	;
				14'b10101001111110: Data_out <= 16'h9244	;
				14'b10101001111111: Data_out <= 16'h923D	;
				14'b10101010000000: Data_out <= 16'h9237	;
				14'b10101010000001: Data_out <= 16'h9230	;
				14'b10101010000010: Data_out <= 16'h922A	;
				14'b10101010000011: Data_out <= 16'h9224	;
				14'b10101010000100: Data_out <= 16'h921D	;
				14'b10101010000101: Data_out <= 16'h9217	;
				14'b10101010000110: Data_out <= 16'h9210	;
				14'b10101010000111: Data_out <= 16'h920A	;
				14'b10101010001000: Data_out <= 16'h9203	;
				14'b10101010001001: Data_out <= 16'h91FD	;
				14'b10101010001010: Data_out <= 16'h91F7	;
				14'b10101010001011: Data_out <= 16'h91F0	;
				14'b10101010001100: Data_out <= 16'h91EA	;
				14'b10101010001101: Data_out <= 16'h91E3	;
				14'b10101010001110: Data_out <= 16'h91DD	;
				14'b10101010001111: Data_out <= 16'h91D6	;
				14'b10101010010000: Data_out <= 16'h91D0	;
				14'b10101010010001: Data_out <= 16'h91CA	;
				14'b10101010010010: Data_out <= 16'h91C3	;
				14'b10101010010011: Data_out <= 16'h91BD	;
				14'b10101010010100: Data_out <= 16'h91B7	;
				14'b10101010010101: Data_out <= 16'h91B0	;
				14'b10101010010110: Data_out <= 16'h91AA	;
				14'b10101010010111: Data_out <= 16'h91A3	;
				14'b10101010011000: Data_out <= 16'h919D	;
				14'b10101010011001: Data_out <= 16'h9197	;
				14'b10101010011010: Data_out <= 16'h9190	;
				14'b10101010011011: Data_out <= 16'h918A	;
				14'b10101010011100: Data_out <= 16'h9184	;
				14'b10101010011101: Data_out <= 16'h917D	;
				14'b10101010011110: Data_out <= 16'h9177	;
				14'b10101010011111: Data_out <= 16'h9171	;
				14'b10101010100000: Data_out <= 16'h916A	;
				14'b10101010100001: Data_out <= 16'h9164	;
				14'b10101010100010: Data_out <= 16'h915E	;
				14'b10101010100011: Data_out <= 16'h9157	;
				14'b10101010100100: Data_out <= 16'h9151	;
				14'b10101010100101: Data_out <= 16'h914B	;
				14'b10101010100110: Data_out <= 16'h9144	;
				14'b10101010100111: Data_out <= 16'h913E	;
				14'b10101010101000: Data_out <= 16'h9138	;
				14'b10101010101001: Data_out <= 16'h9132	;
				14'b10101010101010: Data_out <= 16'h912B	;
				14'b10101010101011: Data_out <= 16'h9125	;
				14'b10101010101100: Data_out <= 16'h911F	;
				14'b10101010101101: Data_out <= 16'h9118	;
				14'b10101010101110: Data_out <= 16'h9112	;
				14'b10101010101111: Data_out <= 16'h910C	;
				14'b10101010110000: Data_out <= 16'h9106	;
				14'b10101010110001: Data_out <= 16'h90FF	;
				14'b10101010110010: Data_out <= 16'h90F9	;
				14'b10101010110011: Data_out <= 16'h90F3	;
				14'b10101010110100: Data_out <= 16'h90ED	;
				14'b10101010110101: Data_out <= 16'h90E6	;
				14'b10101010110110: Data_out <= 16'h90E0	;
				14'b10101010110111: Data_out <= 16'h90DA	;
				14'b10101010111000: Data_out <= 16'h90D4	;
				14'b10101010111001: Data_out <= 16'h90CD	;
				14'b10101010111010: Data_out <= 16'h90C7	;
				14'b10101010111011: Data_out <= 16'h90C1	;
				14'b10101010111100: Data_out <= 16'h90BB	;
				14'b10101010111101: Data_out <= 16'h90B5	;
				14'b10101010111110: Data_out <= 16'h90AE	;
				14'b10101010111111: Data_out <= 16'h90A8	;
				14'b10101011000000: Data_out <= 16'h90A2	;
				14'b10101011000001: Data_out <= 16'h909C	;
				14'b10101011000010: Data_out <= 16'h9096	;
				14'b10101011000011: Data_out <= 16'h908F	;
				14'b10101011000100: Data_out <= 16'h9089	;
				14'b10101011000101: Data_out <= 16'h9083	;
				14'b10101011000110: Data_out <= 16'h907D	;
				14'b10101011000111: Data_out <= 16'h9077	;
				14'b10101011001000: Data_out <= 16'h9071	;
				14'b10101011001001: Data_out <= 16'h906A	;
				14'b10101011001010: Data_out <= 16'h9064	;
				14'b10101011001011: Data_out <= 16'h905E	;
				14'b10101011001100: Data_out <= 16'h9058	;
				14'b10101011001101: Data_out <= 16'h9052	;
				14'b10101011001110: Data_out <= 16'h904C	;
				14'b10101011001111: Data_out <= 16'h9046	;
				14'b10101011010000: Data_out <= 16'h903F	;
				14'b10101011010001: Data_out <= 16'h9039	;
				14'b10101011010010: Data_out <= 16'h9033	;
				14'b10101011010011: Data_out <= 16'h902D	;
				14'b10101011010100: Data_out <= 16'h9027	;
				14'b10101011010101: Data_out <= 16'h9021	;
				14'b10101011010110: Data_out <= 16'h901B	;
				14'b10101011010111: Data_out <= 16'h9015	;
				14'b10101011011000: Data_out <= 16'h900F	;
				14'b10101011011001: Data_out <= 16'h9008	;
				14'b10101011011010: Data_out <= 16'h9002	;
				14'b10101011011011: Data_out <= 16'h8FFC	;
				14'b10101011011100: Data_out <= 16'h8FF6	;
				14'b10101011011101: Data_out <= 16'h8FF0	;
				14'b10101011011110: Data_out <= 16'h8FEA	;
				14'b10101011011111: Data_out <= 16'h8FE4	;
				14'b10101011100000: Data_out <= 16'h8FDE	;
				14'b10101011100001: Data_out <= 16'h8FD8	;
				14'b10101011100010: Data_out <= 16'h8FD2	;
				14'b10101011100011: Data_out <= 16'h8FCC	;
				14'b10101011100100: Data_out <= 16'h8FC6	;
				14'b10101011100101: Data_out <= 16'h8FC0	;
				14'b10101011100110: Data_out <= 16'h8FBA	;
				14'b10101011100111: Data_out <= 16'h8FB4	;
				14'b10101011101000: Data_out <= 16'h8FAE	;
				14'b10101011101001: Data_out <= 16'h8FA8	;
				14'b10101011101010: Data_out <= 16'h8FA2	;
				14'b10101011101011: Data_out <= 16'h8F9C	;
				14'b10101011101100: Data_out <= 16'h8F96	;
				14'b10101011101101: Data_out <= 16'h8F8F	;
				14'b10101011101110: Data_out <= 16'h8F89	;
				14'b10101011101111: Data_out <= 16'h8F83	;
				14'b10101011110000: Data_out <= 16'h8F7E	;
				14'b10101011110001: Data_out <= 16'h8F78	;
				14'b10101011110010: Data_out <= 16'h8F72	;
				14'b10101011110011: Data_out <= 16'h8F6C	;
				14'b10101011110100: Data_out <= 16'h8F66	;
				14'b10101011110101: Data_out <= 16'h8F60	;
				14'b10101011110110: Data_out <= 16'h8F5A	;
				14'b10101011110111: Data_out <= 16'h8F54	;
				14'b10101011111000: Data_out <= 16'h8F4E	;
				14'b10101011111001: Data_out <= 16'h8F48	;
				14'b10101011111010: Data_out <= 16'h8F42	;
				14'b10101011111011: Data_out <= 16'h8F3C	;
				14'b10101011111100: Data_out <= 16'h8F36	;
				14'b10101011111101: Data_out <= 16'h8F30	;
				14'b10101011111110: Data_out <= 16'h8F2A	;
				14'b10101011111111: Data_out <= 16'h8F24	;
				14'b10101100000000: Data_out <= 16'h8F1E	;
				14'b10101100000001: Data_out <= 16'h8F18	;
				14'b10101100000010: Data_out <= 16'h8F12	;
				14'b10101100000011: Data_out <= 16'h8F0C	;
				14'b10101100000100: Data_out <= 16'h8F07	;
				14'b10101100000101: Data_out <= 16'h8F01	;
				14'b10101100000110: Data_out <= 16'h8EFB	;
				14'b10101100000111: Data_out <= 16'h8EF5	;
				14'b10101100001000: Data_out <= 16'h8EEF	;
				14'b10101100001001: Data_out <= 16'h8EE9	;
				14'b10101100001010: Data_out <= 16'h8EE3	;
				14'b10101100001011: Data_out <= 16'h8EDD	;
				14'b10101100001100: Data_out <= 16'h8ED7	;
				14'b10101100001101: Data_out <= 16'h8ED2	;
				14'b10101100001110: Data_out <= 16'h8ECC	;
				14'b10101100001111: Data_out <= 16'h8EC6	;
				14'b10101100010000: Data_out <= 16'h8EC0	;
				14'b10101100010001: Data_out <= 16'h8EBA	;
				14'b10101100010010: Data_out <= 16'h8EB4	;
				14'b10101100010011: Data_out <= 16'h8EAE	;
				14'b10101100010100: Data_out <= 16'h8EA9	;
				14'b10101100010101: Data_out <= 16'h8EA3	;
				14'b10101100010110: Data_out <= 16'h8E9D	;
				14'b10101100010111: Data_out <= 16'h8E97	;
				14'b10101100011000: Data_out <= 16'h8E91	;
				14'b10101100011001: Data_out <= 16'h8E8B	;
				14'b10101100011010: Data_out <= 16'h8E86	;
				14'b10101100011011: Data_out <= 16'h8E80	;
				14'b10101100011100: Data_out <= 16'h8E7A	;
				14'b10101100011101: Data_out <= 16'h8E74	;
				14'b10101100011110: Data_out <= 16'h8E6E	;
				14'b10101100011111: Data_out <= 16'h8E69	;
				14'b10101100100000: Data_out <= 16'h8E63	;
				14'b10101100100001: Data_out <= 16'h8E5D	;
				14'b10101100100010: Data_out <= 16'h8E57	;
				14'b10101100100011: Data_out <= 16'h8E51	;
				14'b10101100100100: Data_out <= 16'h8E4C	;
				14'b10101100100101: Data_out <= 16'h8E46	;
				14'b10101100100110: Data_out <= 16'h8E40	;
				14'b10101100100111: Data_out <= 16'h8E3A	;
				14'b10101100101000: Data_out <= 16'h8E35	;
				14'b10101100101001: Data_out <= 16'h8E2F	;
				14'b10101100101010: Data_out <= 16'h8E29	;
				14'b10101100101011: Data_out <= 16'h8E23	;
				14'b10101100101100: Data_out <= 16'h8E1E	;
				14'b10101100101101: Data_out <= 16'h8E18	;
				14'b10101100101110: Data_out <= 16'h8E12	;
				14'b10101100101111: Data_out <= 16'h8E0C	;
				14'b10101100110000: Data_out <= 16'h8E07	;
				14'b10101100110001: Data_out <= 16'h8E01	;
				14'b10101100110010: Data_out <= 16'h8DFB	;
				14'b10101100110011: Data_out <= 16'h8DF6	;
				14'b10101100110100: Data_out <= 16'h8DF0	;
				14'b10101100110101: Data_out <= 16'h8DEA	;
				14'b10101100110110: Data_out <= 16'h8DE5	;
				14'b10101100110111: Data_out <= 16'h8DDF	;
				14'b10101100111000: Data_out <= 16'h8DD9	;
				14'b10101100111001: Data_out <= 16'h8DD3	;
				14'b10101100111010: Data_out <= 16'h8DCE	;
				14'b10101100111011: Data_out <= 16'h8DC8	;
				14'b10101100111100: Data_out <= 16'h8DC2	;
				14'b10101100111101: Data_out <= 16'h8DBD	;
				14'b10101100111110: Data_out <= 16'h8DB7	;
				14'b10101100111111: Data_out <= 16'h8DB1	;
				14'b10101101000000: Data_out <= 16'h8DAC	;
				14'b10101101000001: Data_out <= 16'h8DA6	;
				14'b10101101000010: Data_out <= 16'h8DA1	;
				14'b10101101000011: Data_out <= 16'h8D9B	;
				14'b10101101000100: Data_out <= 16'h8D95	;
				14'b10101101000101: Data_out <= 16'h8D90	;
				14'b10101101000110: Data_out <= 16'h8D8A	;
				14'b10101101000111: Data_out <= 16'h8D84	;
				14'b10101101001000: Data_out <= 16'h8D7F	;
				14'b10101101001001: Data_out <= 16'h8D79	;
				14'b10101101001010: Data_out <= 16'h8D74	;
				14'b10101101001011: Data_out <= 16'h8D6E	;
				14'b10101101001100: Data_out <= 16'h8D68	;
				14'b10101101001101: Data_out <= 16'h8D63	;
				14'b10101101001110: Data_out <= 16'h8D5D	;
				14'b10101101001111: Data_out <= 16'h8D58	;
				14'b10101101010000: Data_out <= 16'h8D52	;
				14'b10101101010001: Data_out <= 16'h8D4C	;
				14'b10101101010010: Data_out <= 16'h8D47	;
				14'b10101101010011: Data_out <= 16'h8D41	;
				14'b10101101010100: Data_out <= 16'h8D3C	;
				14'b10101101010101: Data_out <= 16'h8D36	;
				14'b10101101010110: Data_out <= 16'h8D31	;
				14'b10101101010111: Data_out <= 16'h8D2B	;
				14'b10101101011000: Data_out <= 16'h8D25	;
				14'b10101101011001: Data_out <= 16'h8D20	;
				14'b10101101011010: Data_out <= 16'h8D1A	;
				14'b10101101011011: Data_out <= 16'h8D15	;
				14'b10101101011100: Data_out <= 16'h8D0F	;
				14'b10101101011101: Data_out <= 16'h8D0A	;
				14'b10101101011110: Data_out <= 16'h8D04	;
				14'b10101101011111: Data_out <= 16'h8CFF	;
				14'b10101101100000: Data_out <= 16'h8CF9	;
				14'b10101101100001: Data_out <= 16'h8CF4	;
				14'b10101101100010: Data_out <= 16'h8CEE	;
				14'b10101101100011: Data_out <= 16'h8CE9	;
				14'b10101101100100: Data_out <= 16'h8CE3	;
				14'b10101101100101: Data_out <= 16'h8CDE	;
				14'b10101101100110: Data_out <= 16'h8CD8	;
				14'b10101101100111: Data_out <= 16'h8CD3	;
				14'b10101101101000: Data_out <= 16'h8CCD	;
				14'b10101101101001: Data_out <= 16'h8CC8	;
				14'b10101101101010: Data_out <= 16'h8CC2	;
				14'b10101101101011: Data_out <= 16'h8CBD	;
				14'b10101101101100: Data_out <= 16'h8CB7	;
				14'b10101101101101: Data_out <= 16'h8CB2	;
				14'b10101101101110: Data_out <= 16'h8CAC	;
				14'b10101101101111: Data_out <= 16'h8CA7	;
				14'b10101101110000: Data_out <= 16'h8CA2	;
				14'b10101101110001: Data_out <= 16'h8C9C	;
				14'b10101101110010: Data_out <= 16'h8C97	;
				14'b10101101110011: Data_out <= 16'h8C91	;
				14'b10101101110100: Data_out <= 16'h8C8C	;
				14'b10101101110101: Data_out <= 16'h8C86	;
				14'b10101101110110: Data_out <= 16'h8C81	;
				14'b10101101110111: Data_out <= 16'h8C7C	;
				14'b10101101111000: Data_out <= 16'h8C76	;
				14'b10101101111001: Data_out <= 16'h8C71	;
				14'b10101101111010: Data_out <= 16'h8C6B	;
				14'b10101101111011: Data_out <= 16'h8C66	;
				14'b10101101111100: Data_out <= 16'h8C61	;
				14'b10101101111101: Data_out <= 16'h8C5B	;
				14'b10101101111110: Data_out <= 16'h8C56	;
				14'b10101101111111: Data_out <= 16'h8C50	;
				14'b10101110000000: Data_out <= 16'h8C4B	;
				14'b10101110000001: Data_out <= 16'h8C46	;
				14'b10101110000010: Data_out <= 16'h8C40	;
				14'b10101110000011: Data_out <= 16'h8C3B	;
				14'b10101110000100: Data_out <= 16'h8C36	;
				14'b10101110000101: Data_out <= 16'h8C30	;
				14'b10101110000110: Data_out <= 16'h8C2B	;
				14'b10101110000111: Data_out <= 16'h8C26	;
				14'b10101110001000: Data_out <= 16'h8C20	;
				14'b10101110001001: Data_out <= 16'h8C1B	;
				14'b10101110001010: Data_out <= 16'h8C16	;
				14'b10101110001011: Data_out <= 16'h8C10	;
				14'b10101110001100: Data_out <= 16'h8C0B	;
				14'b10101110001101: Data_out <= 16'h8C06	;
				14'b10101110001110: Data_out <= 16'h8C00	;
				14'b10101110001111: Data_out <= 16'h8BFB	;
				14'b10101110010000: Data_out <= 16'h8BF6	;
				14'b10101110010001: Data_out <= 16'h8BF0	;
				14'b10101110010010: Data_out <= 16'h8BEB	;
				14'b10101110010011: Data_out <= 16'h8BE6	;
				14'b10101110010100: Data_out <= 16'h8BE1	;
				14'b10101110010101: Data_out <= 16'h8BDB	;
				14'b10101110010110: Data_out <= 16'h8BD6	;
				14'b10101110010111: Data_out <= 16'h8BD1	;
				14'b10101110011000: Data_out <= 16'h8BCB	;
				14'b10101110011001: Data_out <= 16'h8BC6	;
				14'b10101110011010: Data_out <= 16'h8BC1	;
				14'b10101110011011: Data_out <= 16'h8BBC	;
				14'b10101110011100: Data_out <= 16'h8BB6	;
				14'b10101110011101: Data_out <= 16'h8BB1	;
				14'b10101110011110: Data_out <= 16'h8BAC	;
				14'b10101110011111: Data_out <= 16'h8BA7	;
				14'b10101110100000: Data_out <= 16'h8BA1	;
				14'b10101110100001: Data_out <= 16'h8B9C	;
				14'b10101110100010: Data_out <= 16'h8B97	;
				14'b10101110100011: Data_out <= 16'h8B92	;
				14'b10101110100100: Data_out <= 16'h8B8C	;
				14'b10101110100101: Data_out <= 16'h8B87	;
				14'b10101110100110: Data_out <= 16'h8B82	;
				14'b10101110100111: Data_out <= 16'h8B7D	;
				14'b10101110101000: Data_out <= 16'h8B78	;
				14'b10101110101001: Data_out <= 16'h8B72	;
				14'b10101110101010: Data_out <= 16'h8B6D	;
				14'b10101110101011: Data_out <= 16'h8B68	;
				14'b10101110101100: Data_out <= 16'h8B63	;
				14'b10101110101101: Data_out <= 16'h8B5E	;
				14'b10101110101110: Data_out <= 16'h8B59	;
				14'b10101110101111: Data_out <= 16'h8B53	;
				14'b10101110110000: Data_out <= 16'h8B4E	;
				14'b10101110110001: Data_out <= 16'h8B49	;
				14'b10101110110010: Data_out <= 16'h8B44	;
				14'b10101110110011: Data_out <= 16'h8B3F	;
				14'b10101110110100: Data_out <= 16'h8B3A	;
				14'b10101110110101: Data_out <= 16'h8B34	;
				14'b10101110110110: Data_out <= 16'h8B2F	;
				14'b10101110110111: Data_out <= 16'h8B2A	;
				14'b10101110111000: Data_out <= 16'h8B25	;
				14'b10101110111001: Data_out <= 16'h8B20	;
				14'b10101110111010: Data_out <= 16'h8B1B	;
				14'b10101110111011: Data_out <= 16'h8B16	;
				14'b10101110111100: Data_out <= 16'h8B11	;
				14'b10101110111101: Data_out <= 16'h8B0B	;
				14'b10101110111110: Data_out <= 16'h8B06	;
				14'b10101110111111: Data_out <= 16'h8B01	;
				14'b10101111000000: Data_out <= 16'h8AFC	;
				14'b10101111000001: Data_out <= 16'h8AF7	;
				14'b10101111000010: Data_out <= 16'h8AF2	;
				14'b10101111000011: Data_out <= 16'h8AED	;
				14'b10101111000100: Data_out <= 16'h8AE8	;
				14'b10101111000101: Data_out <= 16'h8AE3	;
				14'b10101111000110: Data_out <= 16'h8ADE	;
				14'b10101111000111: Data_out <= 16'h8AD9	;
				14'b10101111001000: Data_out <= 16'h8AD4	;
				14'b10101111001001: Data_out <= 16'h8ACF	;
				14'b10101111001010: Data_out <= 16'h8AC9	;
				14'b10101111001011: Data_out <= 16'h8AC4	;
				14'b10101111001100: Data_out <= 16'h8ABF	;
				14'b10101111001101: Data_out <= 16'h8ABA	;
				14'b10101111001110: Data_out <= 16'h8AB5	;
				14'b10101111001111: Data_out <= 16'h8AB0	;
				14'b10101111010000: Data_out <= 16'h8AAB	;
				14'b10101111010001: Data_out <= 16'h8AA6	;
				14'b10101111010010: Data_out <= 16'h8AA1	;
				14'b10101111010011: Data_out <= 16'h8A9C	;
				14'b10101111010100: Data_out <= 16'h8A97	;
				14'b10101111010101: Data_out <= 16'h8A92	;
				14'b10101111010110: Data_out <= 16'h8A8D	;
				14'b10101111010111: Data_out <= 16'h8A88	;
				14'b10101111011000: Data_out <= 16'h8A83	;
				14'b10101111011001: Data_out <= 16'h8A7E	;
				14'b10101111011010: Data_out <= 16'h8A79	;
				14'b10101111011011: Data_out <= 16'h8A74	;
				14'b10101111011100: Data_out <= 16'h8A6F	;
				14'b10101111011101: Data_out <= 16'h8A6A	;
				14'b10101111011110: Data_out <= 16'h8A65	;
				14'b10101111011111: Data_out <= 16'h8A60	;
				14'b10101111100000: Data_out <= 16'h8A5B	;
				14'b10101111100001: Data_out <= 16'h8A57	;
				14'b10101111100010: Data_out <= 16'h8A52	;
				14'b10101111100011: Data_out <= 16'h8A4D	;
				14'b10101111100100: Data_out <= 16'h8A48	;
				14'b10101111100101: Data_out <= 16'h8A43	;
				14'b10101111100110: Data_out <= 16'h8A3E	;
				14'b10101111100111: Data_out <= 16'h8A39	;
				14'b10101111101000: Data_out <= 16'h8A34	;
				14'b10101111101001: Data_out <= 16'h8A2F	;
				14'b10101111101010: Data_out <= 16'h8A2A	;
				14'b10101111101011: Data_out <= 16'h8A25	;
				14'b10101111101100: Data_out <= 16'h8A20	;
				14'b10101111101101: Data_out <= 16'h8A1C	;
				14'b10101111101110: Data_out <= 16'h8A17	;
				14'b10101111101111: Data_out <= 16'h8A12	;
				14'b10101111110000: Data_out <= 16'h8A0D	;
				14'b10101111110001: Data_out <= 16'h8A08	;
				14'b10101111110010: Data_out <= 16'h8A03	;
				14'b10101111110011: Data_out <= 16'h89FE	;
				14'b10101111110100: Data_out <= 16'h89F9	;
				14'b10101111110101: Data_out <= 16'h89F5	;
				14'b10101111110110: Data_out <= 16'h89F0	;
				14'b10101111110111: Data_out <= 16'h89EB	;
				14'b10101111111000: Data_out <= 16'h89E6	;
				14'b10101111111001: Data_out <= 16'h89E1	;
				14'b10101111111010: Data_out <= 16'h89DC	;
				14'b10101111111011: Data_out <= 16'h89D7	;
				14'b10101111111100: Data_out <= 16'h89D3	;
				14'b10101111111101: Data_out <= 16'h89CE	;
				14'b10101111111110: Data_out <= 16'h89C9	;
				14'b10101111111111: Data_out <= 16'h89C4	;
				14'b10110000000000: Data_out <= 16'h89BF	;
				14'b10110000000001: Data_out <= 16'h89BB	;
				14'b10110000000010: Data_out <= 16'h89B6	;
				14'b10110000000011: Data_out <= 16'h89B1	;
				14'b10110000000100: Data_out <= 16'h89AC	;
				14'b10110000000101: Data_out <= 16'h89A7	;
				14'b10110000000110: Data_out <= 16'h89A3	;
				14'b10110000000111: Data_out <= 16'h899E	;
				14'b10110000001000: Data_out <= 16'h8999	;
				14'b10110000001001: Data_out <= 16'h8994	;
				14'b10110000001010: Data_out <= 16'h898F	;
				14'b10110000001011: Data_out <= 16'h898B	;
				14'b10110000001100: Data_out <= 16'h8986	;
				14'b10110000001101: Data_out <= 16'h8981	;
				14'b10110000001110: Data_out <= 16'h897C	;
				14'b10110000001111: Data_out <= 16'h8978	;
				14'b10110000010000: Data_out <= 16'h8973	;
				14'b10110000010001: Data_out <= 16'h896E	;
				14'b10110000010010: Data_out <= 16'h896A	;
				14'b10110000010011: Data_out <= 16'h8965	;
				14'b10110000010100: Data_out <= 16'h8960	;
				14'b10110000010101: Data_out <= 16'h895B	;
				14'b10110000010110: Data_out <= 16'h8957	;
				14'b10110000010111: Data_out <= 16'h8952	;
				14'b10110000011000: Data_out <= 16'h894D	;
				14'b10110000011001: Data_out <= 16'h8949	;
				14'b10110000011010: Data_out <= 16'h8944	;
				14'b10110000011011: Data_out <= 16'h893F	;
				14'b10110000011100: Data_out <= 16'h893A	;
				14'b10110000011101: Data_out <= 16'h8936	;
				14'b10110000011110: Data_out <= 16'h8931	;
				14'b10110000011111: Data_out <= 16'h892C	;
				14'b10110000100000: Data_out <= 16'h8928	;
				14'b10110000100001: Data_out <= 16'h8923	;
				14'b10110000100010: Data_out <= 16'h891E	;
				14'b10110000100011: Data_out <= 16'h891A	;
				14'b10110000100100: Data_out <= 16'h8915	;
				14'b10110000100101: Data_out <= 16'h8910	;
				14'b10110000100110: Data_out <= 16'h890C	;
				14'b10110000100111: Data_out <= 16'h8907	;
				14'b10110000101000: Data_out <= 16'h8903	;
				14'b10110000101001: Data_out <= 16'h88FE	;
				14'b10110000101010: Data_out <= 16'h88F9	;
				14'b10110000101011: Data_out <= 16'h88F5	;
				14'b10110000101100: Data_out <= 16'h88F0	;
				14'b10110000101101: Data_out <= 16'h88EB	;
				14'b10110000101110: Data_out <= 16'h88E7	;
				14'b10110000101111: Data_out <= 16'h88E2	;
				14'b10110000110000: Data_out <= 16'h88DE	;
				14'b10110000110001: Data_out <= 16'h88D9	;
				14'b10110000110010: Data_out <= 16'h88D4	;
				14'b10110000110011: Data_out <= 16'h88D0	;
				14'b10110000110100: Data_out <= 16'h88CB	;
				14'b10110000110101: Data_out <= 16'h88C7	;
				14'b10110000110110: Data_out <= 16'h88C2	;
				14'b10110000110111: Data_out <= 16'h88BE	;
				14'b10110000111000: Data_out <= 16'h88B9	;
				14'b10110000111001: Data_out <= 16'h88B4	;
				14'b10110000111010: Data_out <= 16'h88B0	;
				14'b10110000111011: Data_out <= 16'h88AB	;
				14'b10110000111100: Data_out <= 16'h88A7	;
				14'b10110000111101: Data_out <= 16'h88A2	;
				14'b10110000111110: Data_out <= 16'h889E	;
				14'b10110000111111: Data_out <= 16'h8899	;
				14'b10110001000000: Data_out <= 16'h8895	;
				14'b10110001000001: Data_out <= 16'h8890	;
				14'b10110001000010: Data_out <= 16'h888C	;
				14'b10110001000011: Data_out <= 16'h8887	;
				14'b10110001000100: Data_out <= 16'h8883	;
				14'b10110001000101: Data_out <= 16'h887E	;
				14'b10110001000110: Data_out <= 16'h887A	;
				14'b10110001000111: Data_out <= 16'h8875	;
				14'b10110001001000: Data_out <= 16'h8871	;
				14'b10110001001001: Data_out <= 16'h886C	;
				14'b10110001001010: Data_out <= 16'h8868	;
				14'b10110001001011: Data_out <= 16'h8863	;
				14'b10110001001100: Data_out <= 16'h885F	;
				14'b10110001001101: Data_out <= 16'h885A	;
				14'b10110001001110: Data_out <= 16'h8856	;
				14'b10110001001111: Data_out <= 16'h8851	;
				14'b10110001010000: Data_out <= 16'h884D	;
				14'b10110001010001: Data_out <= 16'h8848	;
				14'b10110001010010: Data_out <= 16'h8844	;
				14'b10110001010011: Data_out <= 16'h8840	;
				14'b10110001010100: Data_out <= 16'h883B	;
				14'b10110001010101: Data_out <= 16'h8837	;
				14'b10110001010110: Data_out <= 16'h8832	;
				14'b10110001010111: Data_out <= 16'h882E	;
				14'b10110001011000: Data_out <= 16'h8829	;
				14'b10110001011001: Data_out <= 16'h8825	;
				14'b10110001011010: Data_out <= 16'h8821	;
				14'b10110001011011: Data_out <= 16'h881C	;
				14'b10110001011100: Data_out <= 16'h8818	;
				14'b10110001011101: Data_out <= 16'h8813	;
				14'b10110001011110: Data_out <= 16'h880F	;
				14'b10110001011111: Data_out <= 16'h880B	;
				14'b10110001100000: Data_out <= 16'h8806	;
				14'b10110001100001: Data_out <= 16'h8802	;
				14'b10110001100010: Data_out <= 16'h87FE	;
				14'b10110001100011: Data_out <= 16'h87F9	;
				14'b10110001100100: Data_out <= 16'h87F5	;
				14'b10110001100101: Data_out <= 16'h87F0	;
				14'b10110001100110: Data_out <= 16'h87EC	;
				14'b10110001100111: Data_out <= 16'h87E8	;
				14'b10110001101000: Data_out <= 16'h87E3	;
				14'b10110001101001: Data_out <= 16'h87DF	;
				14'b10110001101010: Data_out <= 16'h87DB	;
				14'b10110001101011: Data_out <= 16'h87D6	;
				14'b10110001101100: Data_out <= 16'h87D2	;
				14'b10110001101101: Data_out <= 16'h87CE	;
				14'b10110001101110: Data_out <= 16'h87C9	;
				14'b10110001101111: Data_out <= 16'h87C5	;
				14'b10110001110000: Data_out <= 16'h87C1	;
				14'b10110001110001: Data_out <= 16'h87BD	;
				14'b10110001110010: Data_out <= 16'h87B8	;
				14'b10110001110011: Data_out <= 16'h87B4	;
				14'b10110001110100: Data_out <= 16'h87B0	;
				14'b10110001110101: Data_out <= 16'h87AB	;
				14'b10110001110110: Data_out <= 16'h87A7	;
				14'b10110001110111: Data_out <= 16'h87A3	;
				14'b10110001111000: Data_out <= 16'h879F	;
				14'b10110001111001: Data_out <= 16'h879A	;
				14'b10110001111010: Data_out <= 16'h8796	;
				14'b10110001111011: Data_out <= 16'h8792	;
				14'b10110001111100: Data_out <= 16'h878D	;
				14'b10110001111101: Data_out <= 16'h8789	;
				14'b10110001111110: Data_out <= 16'h8785	;
				14'b10110001111111: Data_out <= 16'h8781	;
				14'b10110010000000: Data_out <= 16'h877D	;
				14'b10110010000001: Data_out <= 16'h8778	;
				14'b10110010000010: Data_out <= 16'h8774	;
				14'b10110010000011: Data_out <= 16'h8770	;
				14'b10110010000100: Data_out <= 16'h876C	;
				14'b10110010000101: Data_out <= 16'h8767	;
				14'b10110010000110: Data_out <= 16'h8763	;
				14'b10110010000111: Data_out <= 16'h875F	;
				14'b10110010001000: Data_out <= 16'h875B	;
				14'b10110010001001: Data_out <= 16'h8757	;
				14'b10110010001010: Data_out <= 16'h8752	;
				14'b10110010001011: Data_out <= 16'h874E	;
				14'b10110010001100: Data_out <= 16'h874A	;
				14'b10110010001101: Data_out <= 16'h8746	;
				14'b10110010001110: Data_out <= 16'h8742	;
				14'b10110010001111: Data_out <= 16'h873E	;
				14'b10110010010000: Data_out <= 16'h8739	;
				14'b10110010010001: Data_out <= 16'h8735	;
				14'b10110010010010: Data_out <= 16'h8731	;
				14'b10110010010011: Data_out <= 16'h872D	;
				14'b10110010010100: Data_out <= 16'h8729	;
				14'b10110010010101: Data_out <= 16'h8725	;
				14'b10110010010110: Data_out <= 16'h8720	;
				14'b10110010010111: Data_out <= 16'h871C	;
				14'b10110010011000: Data_out <= 16'h8718	;
				14'b10110010011001: Data_out <= 16'h8714	;
				14'b10110010011010: Data_out <= 16'h8710	;
				14'b10110010011011: Data_out <= 16'h870C	;
				14'b10110010011100: Data_out <= 16'h8708	;
				14'b10110010011101: Data_out <= 16'h8704	;
				14'b10110010011110: Data_out <= 16'h8700	;
				14'b10110010011111: Data_out <= 16'h86FB	;
				14'b10110010100000: Data_out <= 16'h86F7	;
				14'b10110010100001: Data_out <= 16'h86F3	;
				14'b10110010100010: Data_out <= 16'h86EF	;
				14'b10110010100011: Data_out <= 16'h86EB	;
				14'b10110010100100: Data_out <= 16'h86E7	;
				14'b10110010100101: Data_out <= 16'h86E3	;
				14'b10110010100110: Data_out <= 16'h86DF	;
				14'b10110010100111: Data_out <= 16'h86DB	;
				14'b10110010101000: Data_out <= 16'h86D7	;
				14'b10110010101001: Data_out <= 16'h86D3	;
				14'b10110010101010: Data_out <= 16'h86CF	;
				14'b10110010101011: Data_out <= 16'h86CB	;
				14'b10110010101100: Data_out <= 16'h86C7	;
				14'b10110010101101: Data_out <= 16'h86C3	;
				14'b10110010101110: Data_out <= 16'h86BF	;
				14'b10110010101111: Data_out <= 16'h86BB	;
				14'b10110010110000: Data_out <= 16'h86B7	;
				14'b10110010110001: Data_out <= 16'h86B3	;
				14'b10110010110010: Data_out <= 16'h86AF	;
				14'b10110010110011: Data_out <= 16'h86AB	;
				14'b10110010110100: Data_out <= 16'h86A7	;
				14'b10110010110101: Data_out <= 16'h86A3	;
				14'b10110010110110: Data_out <= 16'h869F	;
				14'b10110010110111: Data_out <= 16'h869B	;
				14'b10110010111000: Data_out <= 16'h8697	;
				14'b10110010111001: Data_out <= 16'h8693	;
				14'b10110010111010: Data_out <= 16'h868F	;
				14'b10110010111011: Data_out <= 16'h868B	;
				14'b10110010111100: Data_out <= 16'h8687	;
				14'b10110010111101: Data_out <= 16'h8683	;
				14'b10110010111110: Data_out <= 16'h867F	;
				14'b10110010111111: Data_out <= 16'h867B	;
				14'b10110011000000: Data_out <= 16'h8677	;
				14'b10110011000001: Data_out <= 16'h8673	;
				14'b10110011000010: Data_out <= 16'h866F	;
				14'b10110011000011: Data_out <= 16'h866B	;
				14'b10110011000100: Data_out <= 16'h8667	;
				14'b10110011000101: Data_out <= 16'h8663	;
				14'b10110011000110: Data_out <= 16'h865F	;
				14'b10110011000111: Data_out <= 16'h865B	;
				14'b10110011001000: Data_out <= 16'h8658	;
				14'b10110011001001: Data_out <= 16'h8654	;
				14'b10110011001010: Data_out <= 16'h8650	;
				14'b10110011001011: Data_out <= 16'h864C	;
				14'b10110011001100: Data_out <= 16'h8648	;
				14'b10110011001101: Data_out <= 16'h8644	;
				14'b10110011001110: Data_out <= 16'h8640	;
				14'b10110011001111: Data_out <= 16'h863C	;
				14'b10110011010000: Data_out <= 16'h8638	;
				14'b10110011010001: Data_out <= 16'h8635	;
				14'b10110011010010: Data_out <= 16'h8631	;
				14'b10110011010011: Data_out <= 16'h862D	;
				14'b10110011010100: Data_out <= 16'h8629	;
				14'b10110011010101: Data_out <= 16'h8625	;
				14'b10110011010110: Data_out <= 16'h8621	;
				14'b10110011010111: Data_out <= 16'h861D	;
				14'b10110011011000: Data_out <= 16'h861A	;
				14'b10110011011001: Data_out <= 16'h8616	;
				14'b10110011011010: Data_out <= 16'h8612	;
				14'b10110011011011: Data_out <= 16'h860E	;
				14'b10110011011100: Data_out <= 16'h860A	;
				14'b10110011011101: Data_out <= 16'h8607	;
				14'b10110011011110: Data_out <= 16'h8603	;
				14'b10110011011111: Data_out <= 16'h85FF	;
				14'b10110011100000: Data_out <= 16'h85FB	;
				14'b10110011100001: Data_out <= 16'h85F7	;
				14'b10110011100010: Data_out <= 16'h85F4	;
				14'b10110011100011: Data_out <= 16'h85F0	;
				14'b10110011100100: Data_out <= 16'h85EC	;
				14'b10110011100101: Data_out <= 16'h85E8	;
				14'b10110011100110: Data_out <= 16'h85E4	;
				14'b10110011100111: Data_out <= 16'h85E1	;
				14'b10110011101000: Data_out <= 16'h85DD	;
				14'b10110011101001: Data_out <= 16'h85D9	;
				14'b10110011101010: Data_out <= 16'h85D5	;
				14'b10110011101011: Data_out <= 16'h85D2	;
				14'b10110011101100: Data_out <= 16'h85CE	;
				14'b10110011101101: Data_out <= 16'h85CA	;
				14'b10110011101110: Data_out <= 16'h85C6	;
				14'b10110011101111: Data_out <= 16'h85C3	;
				14'b10110011110000: Data_out <= 16'h85BF	;
				14'b10110011110001: Data_out <= 16'h85BB	;
				14'b10110011110010: Data_out <= 16'h85B8	;
				14'b10110011110011: Data_out <= 16'h85B4	;
				14'b10110011110100: Data_out <= 16'h85B0	;
				14'b10110011110101: Data_out <= 16'h85AC	;
				14'b10110011110110: Data_out <= 16'h85A9	;
				14'b10110011110111: Data_out <= 16'h85A5	;
				14'b10110011111000: Data_out <= 16'h85A1	;
				14'b10110011111001: Data_out <= 16'h859E	;
				14'b10110011111010: Data_out <= 16'h859A	;
				14'b10110011111011: Data_out <= 16'h8596	;
				14'b10110011111100: Data_out <= 16'h8593	;
				14'b10110011111101: Data_out <= 16'h858F	;
				14'b10110011111110: Data_out <= 16'h858B	;
				14'b10110011111111: Data_out <= 16'h8588	;
				14'b10110100000000: Data_out <= 16'h8584	;
				14'b10110100000001: Data_out <= 16'h8580	;
				14'b10110100000010: Data_out <= 16'h857D	;
				14'b10110100000011: Data_out <= 16'h8579	;
				14'b10110100000100: Data_out <= 16'h8575	;
				14'b10110100000101: Data_out <= 16'h8572	;
				14'b10110100000110: Data_out <= 16'h856E	;
				14'b10110100000111: Data_out <= 16'h856B	;
				14'b10110100001000: Data_out <= 16'h8567	;
				14'b10110100001001: Data_out <= 16'h8563	;
				14'b10110100001010: Data_out <= 16'h8560	;
				14'b10110100001011: Data_out <= 16'h855C	;
				14'b10110100001100: Data_out <= 16'h8559	;
				14'b10110100001101: Data_out <= 16'h8555	;
				14'b10110100001110: Data_out <= 16'h8551	;
				14'b10110100001111: Data_out <= 16'h854E	;
				14'b10110100010000: Data_out <= 16'h854A	;
				14'b10110100010001: Data_out <= 16'h8547	;
				14'b10110100010010: Data_out <= 16'h8543	;
				14'b10110100010011: Data_out <= 16'h8540	;
				14'b10110100010100: Data_out <= 16'h853C	;
				14'b10110100010101: Data_out <= 16'h8538	;
				14'b10110100010110: Data_out <= 16'h8535	;
				14'b10110100010111: Data_out <= 16'h8531	;
				14'b10110100011000: Data_out <= 16'h852E	;
				14'b10110100011001: Data_out <= 16'h852A	;
				14'b10110100011010: Data_out <= 16'h8527	;
				14'b10110100011011: Data_out <= 16'h8523	;
				14'b10110100011100: Data_out <= 16'h8520	;
				14'b10110100011101: Data_out <= 16'h851C	;
				14'b10110100011110: Data_out <= 16'h8519	;
				14'b10110100011111: Data_out <= 16'h8515	;
				14'b10110100100000: Data_out <= 16'h8512	;
				14'b10110100100001: Data_out <= 16'h850E	;
				14'b10110100100010: Data_out <= 16'h850B	;
				14'b10110100100011: Data_out <= 16'h8507	;
				14'b10110100100100: Data_out <= 16'h8504	;
				14'b10110100100101: Data_out <= 16'h8500	;
				14'b10110100100110: Data_out <= 16'h84FD	;
				14'b10110100100111: Data_out <= 16'h84F9	;
				14'b10110100101000: Data_out <= 16'h84F6	;
				14'b10110100101001: Data_out <= 16'h84F2	;
				14'b10110100101010: Data_out <= 16'h84EF	;
				14'b10110100101011: Data_out <= 16'h84EB	;
				14'b10110100101100: Data_out <= 16'h84E8	;
				14'b10110100101101: Data_out <= 16'h84E5	;
				14'b10110100101110: Data_out <= 16'h84E1	;
				14'b10110100101111: Data_out <= 16'h84DE	;
				14'b10110100110000: Data_out <= 16'h84DA	;
				14'b10110100110001: Data_out <= 16'h84D7	;
				14'b10110100110010: Data_out <= 16'h84D3	;
				14'b10110100110011: Data_out <= 16'h84D0	;
				14'b10110100110100: Data_out <= 16'h84CD	;
				14'b10110100110101: Data_out <= 16'h84C9	;
				14'b10110100110110: Data_out <= 16'h84C6	;
				14'b10110100110111: Data_out <= 16'h84C2	;
				14'b10110100111000: Data_out <= 16'h84BF	;
				14'b10110100111001: Data_out <= 16'h84BC	;
				14'b10110100111010: Data_out <= 16'h84B8	;
				14'b10110100111011: Data_out <= 16'h84B5	;
				14'b10110100111100: Data_out <= 16'h84B1	;
				14'b10110100111101: Data_out <= 16'h84AE	;
				14'b10110100111110: Data_out <= 16'h84AB	;
				14'b10110100111111: Data_out <= 16'h84A7	;
				14'b10110101000000: Data_out <= 16'h84A4	;
				14'b10110101000001: Data_out <= 16'h84A1	;
				14'b10110101000010: Data_out <= 16'h849D	;
				14'b10110101000011: Data_out <= 16'h849A	;
				14'b10110101000100: Data_out <= 16'h8497	;
				14'b10110101000101: Data_out <= 16'h8493	;
				14'b10110101000110: Data_out <= 16'h8490	;
				14'b10110101000111: Data_out <= 16'h848D	;
				14'b10110101001000: Data_out <= 16'h8489	;
				14'b10110101001001: Data_out <= 16'h8486	;
				14'b10110101001010: Data_out <= 16'h8483	;
				14'b10110101001011: Data_out <= 16'h847F	;
				14'b10110101001100: Data_out <= 16'h847C	;
				14'b10110101001101: Data_out <= 16'h8479	;
				14'b10110101001110: Data_out <= 16'h8476	;
				14'b10110101001111: Data_out <= 16'h8472	;
				14'b10110101010000: Data_out <= 16'h846F	;
				14'b10110101010001: Data_out <= 16'h846C	;
				14'b10110101010010: Data_out <= 16'h8468	;
				14'b10110101010011: Data_out <= 16'h8465	;
				14'b10110101010100: Data_out <= 16'h8462	;
				14'b10110101010101: Data_out <= 16'h845F	;
				14'b10110101010110: Data_out <= 16'h845B	;
				14'b10110101010111: Data_out <= 16'h8458	;
				14'b10110101011000: Data_out <= 16'h8455	;
				14'b10110101011001: Data_out <= 16'h8452	;
				14'b10110101011010: Data_out <= 16'h844E	;
				14'b10110101011011: Data_out <= 16'h844B	;
				14'b10110101011100: Data_out <= 16'h8448	;
				14'b10110101011101: Data_out <= 16'h8445	;
				14'b10110101011110: Data_out <= 16'h8442	;
				14'b10110101011111: Data_out <= 16'h843E	;
				14'b10110101100000: Data_out <= 16'h843B	;
				14'b10110101100001: Data_out <= 16'h8438	;
				14'b10110101100010: Data_out <= 16'h8435	;
				14'b10110101100011: Data_out <= 16'h8432	;
				14'b10110101100100: Data_out <= 16'h842E	;
				14'b10110101100101: Data_out <= 16'h842B	;
				14'b10110101100110: Data_out <= 16'h8428	;
				14'b10110101100111: Data_out <= 16'h8425	;
				14'b10110101101000: Data_out <= 16'h8422	;
				14'b10110101101001: Data_out <= 16'h841F	;
				14'b10110101101010: Data_out <= 16'h841B	;
				14'b10110101101011: Data_out <= 16'h8418	;
				14'b10110101101100: Data_out <= 16'h8415	;
				14'b10110101101101: Data_out <= 16'h8412	;
				14'b10110101101110: Data_out <= 16'h840F	;
				14'b10110101101111: Data_out <= 16'h840C	;
				14'b10110101110000: Data_out <= 16'h8409	;
				14'b10110101110001: Data_out <= 16'h8405	;
				14'b10110101110010: Data_out <= 16'h8402	;
				14'b10110101110011: Data_out <= 16'h83FF	;
				14'b10110101110100: Data_out <= 16'h83FC	;
				14'b10110101110101: Data_out <= 16'h83F9	;
				14'b10110101110110: Data_out <= 16'h83F6	;
				14'b10110101110111: Data_out <= 16'h83F3	;
				14'b10110101111000: Data_out <= 16'h83F0	;
				14'b10110101111001: Data_out <= 16'h83ED	;
				14'b10110101111010: Data_out <= 16'h83E9	;
				14'b10110101111011: Data_out <= 16'h83E6	;
				14'b10110101111100: Data_out <= 16'h83E3	;
				14'b10110101111101: Data_out <= 16'h83E0	;
				14'b10110101111110: Data_out <= 16'h83DD	;
				14'b10110101111111: Data_out <= 16'h83DA	;
				14'b10110110000000: Data_out <= 16'h83D7	;
				14'b10110110000001: Data_out <= 16'h83D4	;
				14'b10110110000010: Data_out <= 16'h83D1	;
				14'b10110110000011: Data_out <= 16'h83CE	;
				14'b10110110000100: Data_out <= 16'h83CB	;
				14'b10110110000101: Data_out <= 16'h83C8	;
				14'b10110110000110: Data_out <= 16'h83C5	;
				14'b10110110000111: Data_out <= 16'h83C2	;
				14'b10110110001000: Data_out <= 16'h83BF	;
				14'b10110110001001: Data_out <= 16'h83BC	;
				14'b10110110001010: Data_out <= 16'h83B9	;
				14'b10110110001011: Data_out <= 16'h83B6	;
				14'b10110110001100: Data_out <= 16'h83B3	;
				14'b10110110001101: Data_out <= 16'h83B0	;
				14'b10110110001110: Data_out <= 16'h83AD	;
				14'b10110110001111: Data_out <= 16'h83AA	;
				14'b10110110010000: Data_out <= 16'h83A7	;
				14'b10110110010001: Data_out <= 16'h83A4	;
				14'b10110110010010: Data_out <= 16'h83A1	;
				14'b10110110010011: Data_out <= 16'h839E	;
				14'b10110110010100: Data_out <= 16'h839B	;
				14'b10110110010101: Data_out <= 16'h8398	;
				14'b10110110010110: Data_out <= 16'h8395	;
				14'b10110110010111: Data_out <= 16'h8392	;
				14'b10110110011000: Data_out <= 16'h838F	;
				14'b10110110011001: Data_out <= 16'h838C	;
				14'b10110110011010: Data_out <= 16'h8389	;
				14'b10110110011011: Data_out <= 16'h8386	;
				14'b10110110011100: Data_out <= 16'h8383	;
				14'b10110110011101: Data_out <= 16'h8381	;
				14'b10110110011110: Data_out <= 16'h837E	;
				14'b10110110011111: Data_out <= 16'h837B	;
				14'b10110110100000: Data_out <= 16'h8378	;
				14'b10110110100001: Data_out <= 16'h8375	;
				14'b10110110100010: Data_out <= 16'h8372	;
				14'b10110110100011: Data_out <= 16'h836F	;
				14'b10110110100100: Data_out <= 16'h836C	;
				14'b10110110100101: Data_out <= 16'h8369	;
				14'b10110110100110: Data_out <= 16'h8366	;
				14'b10110110100111: Data_out <= 16'h8364	;
				14'b10110110101000: Data_out <= 16'h8361	;
				14'b10110110101001: Data_out <= 16'h835E	;
				14'b10110110101010: Data_out <= 16'h835B	;
				14'b10110110101011: Data_out <= 16'h8358	;
				14'b10110110101100: Data_out <= 16'h8355	;
				14'b10110110101101: Data_out <= 16'h8352	;
				14'b10110110101110: Data_out <= 16'h8350	;
				14'b10110110101111: Data_out <= 16'h834D	;
				14'b10110110110000: Data_out <= 16'h834A	;
				14'b10110110110001: Data_out <= 16'h8347	;
				14'b10110110110010: Data_out <= 16'h8344	;
				14'b10110110110011: Data_out <= 16'h8341	;
				14'b10110110110100: Data_out <= 16'h833F	;
				14'b10110110110101: Data_out <= 16'h833C	;
				14'b10110110110110: Data_out <= 16'h8339	;
				14'b10110110110111: Data_out <= 16'h8336	;
				14'b10110110111000: Data_out <= 16'h8333	;
				14'b10110110111001: Data_out <= 16'h8331	;
				14'b10110110111010: Data_out <= 16'h832E	;
				14'b10110110111011: Data_out <= 16'h832B	;
				14'b10110110111100: Data_out <= 16'h8328	;
				14'b10110110111101: Data_out <= 16'h8326	;
				14'b10110110111110: Data_out <= 16'h8323	;
				14'b10110110111111: Data_out <= 16'h8320	;
				14'b10110111000000: Data_out <= 16'h831D	;
				14'b10110111000001: Data_out <= 16'h831B	;
				14'b10110111000010: Data_out <= 16'h8318	;
				14'b10110111000011: Data_out <= 16'h8315	;
				14'b10110111000100: Data_out <= 16'h8312	;
				14'b10110111000101: Data_out <= 16'h8310	;
				14'b10110111000110: Data_out <= 16'h830D	;
				14'b10110111000111: Data_out <= 16'h830A	;
				14'b10110111001000: Data_out <= 16'h8307	;
				14'b10110111001001: Data_out <= 16'h8305	;
				14'b10110111001010: Data_out <= 16'h8302	;
				14'b10110111001011: Data_out <= 16'h82FF	;
				14'b10110111001100: Data_out <= 16'h82FD	;
				14'b10110111001101: Data_out <= 16'h82FA	;
				14'b10110111001110: Data_out <= 16'h82F7	;
				14'b10110111001111: Data_out <= 16'h82F4	;
				14'b10110111010000: Data_out <= 16'h82F2	;
				14'b10110111010001: Data_out <= 16'h82EF	;
				14'b10110111010010: Data_out <= 16'h82EC	;
				14'b10110111010011: Data_out <= 16'h82EA	;
				14'b10110111010100: Data_out <= 16'h82E7	;
				14'b10110111010101: Data_out <= 16'h82E4	;
				14'b10110111010110: Data_out <= 16'h82E2	;
				14'b10110111010111: Data_out <= 16'h82DF	;
				14'b10110111011000: Data_out <= 16'h82DD	;
				14'b10110111011001: Data_out <= 16'h82DA	;
				14'b10110111011010: Data_out <= 16'h82D7	;
				14'b10110111011011: Data_out <= 16'h82D5	;
				14'b10110111011100: Data_out <= 16'h82D2	;
				14'b10110111011101: Data_out <= 16'h82CF	;
				14'b10110111011110: Data_out <= 16'h82CD	;
				14'b10110111011111: Data_out <= 16'h82CA	;
				14'b10110111100000: Data_out <= 16'h82C8	;
				14'b10110111100001: Data_out <= 16'h82C5	;
				14'b10110111100010: Data_out <= 16'h82C2	;
				14'b10110111100011: Data_out <= 16'h82C0	;
				14'b10110111100100: Data_out <= 16'h82BD	;
				14'b10110111100101: Data_out <= 16'h82BB	;
				14'b10110111100110: Data_out <= 16'h82B8	;
				14'b10110111100111: Data_out <= 16'h82B5	;
				14'b10110111101000: Data_out <= 16'h82B3	;
				14'b10110111101001: Data_out <= 16'h82B0	;
				14'b10110111101010: Data_out <= 16'h82AE	;
				14'b10110111101011: Data_out <= 16'h82AB	;
				14'b10110111101100: Data_out <= 16'h82A9	;
				14'b10110111101101: Data_out <= 16'h82A6	;
				14'b10110111101110: Data_out <= 16'h82A4	;
				14'b10110111101111: Data_out <= 16'h82A1	;
				14'b10110111110000: Data_out <= 16'h829F	;
				14'b10110111110001: Data_out <= 16'h829C	;
				14'b10110111110010: Data_out <= 16'h8299	;
				14'b10110111110011: Data_out <= 16'h8297	;
				14'b10110111110100: Data_out <= 16'h8294	;
				14'b10110111110101: Data_out <= 16'h8292	;
				14'b10110111110110: Data_out <= 16'h828F	;
				14'b10110111110111: Data_out <= 16'h828D	;
				14'b10110111111000: Data_out <= 16'h828A	;
				14'b10110111111001: Data_out <= 16'h8288	;
				14'b10110111111010: Data_out <= 16'h8286	;
				14'b10110111111011: Data_out <= 16'h8283	;
				14'b10110111111100: Data_out <= 16'h8281	;
				14'b10110111111101: Data_out <= 16'h827E	;
				14'b10110111111110: Data_out <= 16'h827C	;
				14'b10110111111111: Data_out <= 16'h8279	;
				14'b10111000000000: Data_out <= 16'h8277	;
				14'b10111000000001: Data_out <= 16'h8274	;
				14'b10111000000010: Data_out <= 16'h8272	;
				14'b10111000000011: Data_out <= 16'h826F	;
				14'b10111000000100: Data_out <= 16'h826D	;
				14'b10111000000101: Data_out <= 16'h826B	;
				14'b10111000000110: Data_out <= 16'h8268	;
				14'b10111000000111: Data_out <= 16'h8266	;
				14'b10111000001000: Data_out <= 16'h8263	;
				14'b10111000001001: Data_out <= 16'h8261	;
				14'b10111000001010: Data_out <= 16'h825E	;
				14'b10111000001011: Data_out <= 16'h825C	;
				14'b10111000001100: Data_out <= 16'h825A	;
				14'b10111000001101: Data_out <= 16'h8257	;
				14'b10111000001110: Data_out <= 16'h8255	;
				14'b10111000001111: Data_out <= 16'h8252	;
				14'b10111000010000: Data_out <= 16'h8250	;
				14'b10111000010001: Data_out <= 16'h824E	;
				14'b10111000010010: Data_out <= 16'h824B	;
				14'b10111000010011: Data_out <= 16'h8249	;
				14'b10111000010100: Data_out <= 16'h8247	;
				14'b10111000010101: Data_out <= 16'h8244	;
				14'b10111000010110: Data_out <= 16'h8242	;
				14'b10111000010111: Data_out <= 16'h8240	;
				14'b10111000011000: Data_out <= 16'h823D	;
				14'b10111000011001: Data_out <= 16'h823B	;
				14'b10111000011010: Data_out <= 16'h8239	;
				14'b10111000011011: Data_out <= 16'h8236	;
				14'b10111000011100: Data_out <= 16'h8234	;
				14'b10111000011101: Data_out <= 16'h8232	;
				14'b10111000011110: Data_out <= 16'h822F	;
				14'b10111000011111: Data_out <= 16'h822D	;
				14'b10111000100000: Data_out <= 16'h822B	;
				14'b10111000100001: Data_out <= 16'h8228	;
				14'b10111000100010: Data_out <= 16'h8226	;
				14'b10111000100011: Data_out <= 16'h8224	;
				14'b10111000100100: Data_out <= 16'h8222	;
				14'b10111000100101: Data_out <= 16'h821F	;
				14'b10111000100110: Data_out <= 16'h821D	;
				14'b10111000100111: Data_out <= 16'h821B	;
				14'b10111000101000: Data_out <= 16'h8218	;
				14'b10111000101001: Data_out <= 16'h8216	;
				14'b10111000101010: Data_out <= 16'h8214	;
				14'b10111000101011: Data_out <= 16'h8212	;
				14'b10111000101100: Data_out <= 16'h820F	;
				14'b10111000101101: Data_out <= 16'h820D	;
				14'b10111000101110: Data_out <= 16'h820B	;
				14'b10111000101111: Data_out <= 16'h8209	;
				14'b10111000110000: Data_out <= 16'h8206	;
				14'b10111000110001: Data_out <= 16'h8204	;
				14'b10111000110010: Data_out <= 16'h8202	;
				14'b10111000110011: Data_out <= 16'h8200	;
				14'b10111000110100: Data_out <= 16'h81FE	;
				14'b10111000110101: Data_out <= 16'h81FB	;
				14'b10111000110110: Data_out <= 16'h81F9	;
				14'b10111000110111: Data_out <= 16'h81F7	;
				14'b10111000111000: Data_out <= 16'h81F5	;
				14'b10111000111001: Data_out <= 16'h81F3	;
				14'b10111000111010: Data_out <= 16'h81F0	;
				14'b10111000111011: Data_out <= 16'h81EE	;
				14'b10111000111100: Data_out <= 16'h81EC	;
				14'b10111000111101: Data_out <= 16'h81EA	;
				14'b10111000111110: Data_out <= 16'h81E8	;
				14'b10111000111111: Data_out <= 16'h81E6	;
				14'b10111001000000: Data_out <= 16'h81E4	;
				14'b10111001000001: Data_out <= 16'h81E1	;
				14'b10111001000010: Data_out <= 16'h81DF	;
				14'b10111001000011: Data_out <= 16'h81DD	;
				14'b10111001000100: Data_out <= 16'h81DB	;
				14'b10111001000101: Data_out <= 16'h81D9	;
				14'b10111001000110: Data_out <= 16'h81D7	;
				14'b10111001000111: Data_out <= 16'h81D5	;
				14'b10111001001000: Data_out <= 16'h81D2	;
				14'b10111001001001: Data_out <= 16'h81D0	;
				14'b10111001001010: Data_out <= 16'h81CE	;
				14'b10111001001011: Data_out <= 16'h81CC	;
				14'b10111001001100: Data_out <= 16'h81CA	;
				14'b10111001001101: Data_out <= 16'h81C8	;
				14'b10111001001110: Data_out <= 16'h81C6	;
				14'b10111001001111: Data_out <= 16'h81C4	;
				14'b10111001010000: Data_out <= 16'h81C2	;
				14'b10111001010001: Data_out <= 16'h81C0	;
				14'b10111001010010: Data_out <= 16'h81BE	;
				14'b10111001010011: Data_out <= 16'h81BC	;
				14'b10111001010100: Data_out <= 16'h81B9	;
				14'b10111001010101: Data_out <= 16'h81B7	;
				14'b10111001010110: Data_out <= 16'h81B5	;
				14'b10111001010111: Data_out <= 16'h81B3	;
				14'b10111001011000: Data_out <= 16'h81B1	;
				14'b10111001011001: Data_out <= 16'h81AF	;
				14'b10111001011010: Data_out <= 16'h81AD	;
				14'b10111001011011: Data_out <= 16'h81AB	;
				14'b10111001011100: Data_out <= 16'h81A9	;
				14'b10111001011101: Data_out <= 16'h81A7	;
				14'b10111001011110: Data_out <= 16'h81A5	;
				14'b10111001011111: Data_out <= 16'h81A3	;
				14'b10111001100000: Data_out <= 16'h81A1	;
				14'b10111001100001: Data_out <= 16'h819F	;
				14'b10111001100010: Data_out <= 16'h819D	;
				14'b10111001100011: Data_out <= 16'h819B	;
				14'b10111001100100: Data_out <= 16'h8199	;
				14'b10111001100101: Data_out <= 16'h8197	;
				14'b10111001100110: Data_out <= 16'h8195	;
				14'b10111001100111: Data_out <= 16'h8193	;
				14'b10111001101000: Data_out <= 16'h8191	;
				14'b10111001101001: Data_out <= 16'h818F	;
				14'b10111001101010: Data_out <= 16'h818D	;
				14'b10111001101011: Data_out <= 16'h818C	;
				14'b10111001101100: Data_out <= 16'h818A	;
				14'b10111001101101: Data_out <= 16'h8188	;
				14'b10111001101110: Data_out <= 16'h8186	;
				14'b10111001101111: Data_out <= 16'h8184	;
				14'b10111001110000: Data_out <= 16'h8182	;
				14'b10111001110001: Data_out <= 16'h8180	;
				14'b10111001110010: Data_out <= 16'h817E	;
				14'b10111001110011: Data_out <= 16'h817C	;
				14'b10111001110100: Data_out <= 16'h817A	;
				14'b10111001110101: Data_out <= 16'h8178	;
				14'b10111001110110: Data_out <= 16'h8176	;
				14'b10111001110111: Data_out <= 16'h8175	;
				14'b10111001111000: Data_out <= 16'h8173	;
				14'b10111001111001: Data_out <= 16'h8171	;
				14'b10111001111010: Data_out <= 16'h816F	;
				14'b10111001111011: Data_out <= 16'h816D	;
				14'b10111001111100: Data_out <= 16'h816B	;
				14'b10111001111101: Data_out <= 16'h8169	;
				14'b10111001111110: Data_out <= 16'h8167	;
				14'b10111001111111: Data_out <= 16'h8166	;
				14'b10111010000000: Data_out <= 16'h8164	;
				14'b10111010000001: Data_out <= 16'h8162	;
				14'b10111010000010: Data_out <= 16'h8160	;
				14'b10111010000011: Data_out <= 16'h815E	;
				14'b10111010000100: Data_out <= 16'h815C	;
				14'b10111010000101: Data_out <= 16'h815B	;
				14'b10111010000110: Data_out <= 16'h8159	;
				14'b10111010000111: Data_out <= 16'h8157	;
				14'b10111010001000: Data_out <= 16'h8155	;
				14'b10111010001001: Data_out <= 16'h8153	;
				14'b10111010001010: Data_out <= 16'h8152	;
				14'b10111010001011: Data_out <= 16'h8150	;
				14'b10111010001100: Data_out <= 16'h814E	;
				14'b10111010001101: Data_out <= 16'h814C	;
				14'b10111010001110: Data_out <= 16'h814A	;
				14'b10111010001111: Data_out <= 16'h8149	;
				14'b10111010010000: Data_out <= 16'h8147	;
				14'b10111010010001: Data_out <= 16'h8145	;
				14'b10111010010010: Data_out <= 16'h8143	;
				14'b10111010010011: Data_out <= 16'h8142	;
				14'b10111010010100: Data_out <= 16'h8140	;
				14'b10111010010101: Data_out <= 16'h813E	;
				14'b10111010010110: Data_out <= 16'h813C	;
				14'b10111010010111: Data_out <= 16'h813B	;
				14'b10111010011000: Data_out <= 16'h8139	;
				14'b10111010011001: Data_out <= 16'h8137	;
				14'b10111010011010: Data_out <= 16'h8135	;
				14'b10111010011011: Data_out <= 16'h8134	;
				14'b10111010011100: Data_out <= 16'h8132	;
				14'b10111010011101: Data_out <= 16'h8130	;
				14'b10111010011110: Data_out <= 16'h812F	;
				14'b10111010011111: Data_out <= 16'h812D	;
				14'b10111010100000: Data_out <= 16'h812B	;
				14'b10111010100001: Data_out <= 16'h812A	;
				14'b10111010100010: Data_out <= 16'h8128	;
				14'b10111010100011: Data_out <= 16'h8126	;
				14'b10111010100100: Data_out <= 16'h8124	;
				14'b10111010100101: Data_out <= 16'h8123	;
				14'b10111010100110: Data_out <= 16'h8121	;
				14'b10111010100111: Data_out <= 16'h811F	;
				14'b10111010101000: Data_out <= 16'h811E	;
				14'b10111010101001: Data_out <= 16'h811C	;
				14'b10111010101010: Data_out <= 16'h811B	;
				14'b10111010101011: Data_out <= 16'h8119	;
				14'b10111010101100: Data_out <= 16'h8117	;
				14'b10111010101101: Data_out <= 16'h8116	;
				14'b10111010101110: Data_out <= 16'h8114	;
				14'b10111010101111: Data_out <= 16'h8112	;
				14'b10111010110000: Data_out <= 16'h8111	;
				14'b10111010110001: Data_out <= 16'h810F	;
				14'b10111010110010: Data_out <= 16'h810E	;
				14'b10111010110011: Data_out <= 16'h810C	;
				14'b10111010110100: Data_out <= 16'h810A	;
				14'b10111010110101: Data_out <= 16'h8109	;
				14'b10111010110110: Data_out <= 16'h8107	;
				14'b10111010110111: Data_out <= 16'h8106	;
				14'b10111010111000: Data_out <= 16'h8104	;
				14'b10111010111001: Data_out <= 16'h8102	;
				14'b10111010111010: Data_out <= 16'h8101	;
				14'b10111010111011: Data_out <= 16'h80FF	;
				14'b10111010111100: Data_out <= 16'h80FE	;
				14'b10111010111101: Data_out <= 16'h80FC	;
				14'b10111010111110: Data_out <= 16'h80FB	;
				14'b10111010111111: Data_out <= 16'h80F9	;
				14'b10111011000000: Data_out <= 16'h80F8	;
				14'b10111011000001: Data_out <= 16'h80F6	;
				14'b10111011000010: Data_out <= 16'h80F4	;
				14'b10111011000011: Data_out <= 16'h80F3	;
				14'b10111011000100: Data_out <= 16'h80F1	;
				14'b10111011000101: Data_out <= 16'h80F0	;
				14'b10111011000110: Data_out <= 16'h80EE	;
				14'b10111011000111: Data_out <= 16'h80ED	;
				14'b10111011001000: Data_out <= 16'h80EB	;
				14'b10111011001001: Data_out <= 16'h80EA	;
				14'b10111011001010: Data_out <= 16'h80E8	;
				14'b10111011001011: Data_out <= 16'h80E7	;
				14'b10111011001100: Data_out <= 16'h80E5	;
				14'b10111011001101: Data_out <= 16'h80E4	;
				14'b10111011001110: Data_out <= 16'h80E2	;
				14'b10111011001111: Data_out <= 16'h80E1	;
				14'b10111011010000: Data_out <= 16'h80E0	;
				14'b10111011010001: Data_out <= 16'h80DE	;
				14'b10111011010010: Data_out <= 16'h80DD	;
				14'b10111011010011: Data_out <= 16'h80DB	;
				14'b10111011010100: Data_out <= 16'h80DA	;
				14'b10111011010101: Data_out <= 16'h80D8	;
				14'b10111011010110: Data_out <= 16'h80D7	;
				14'b10111011010111: Data_out <= 16'h80D5	;
				14'b10111011011000: Data_out <= 16'h80D4	;
				14'b10111011011001: Data_out <= 16'h80D3	;
				14'b10111011011010: Data_out <= 16'h80D1	;
				14'b10111011011011: Data_out <= 16'h80D0	;
				14'b10111011011100: Data_out <= 16'h80CE	;
				14'b10111011011101: Data_out <= 16'h80CD	;
				14'b10111011011110: Data_out <= 16'h80CC	;
				14'b10111011011111: Data_out <= 16'h80CA	;
				14'b10111011100000: Data_out <= 16'h80C9	;
				14'b10111011100001: Data_out <= 16'h80C7	;
				14'b10111011100010: Data_out <= 16'h80C6	;
				14'b10111011100011: Data_out <= 16'h80C5	;
				14'b10111011100100: Data_out <= 16'h80C3	;
				14'b10111011100101: Data_out <= 16'h80C2	;
				14'b10111011100110: Data_out <= 16'h80C1	;
				14'b10111011100111: Data_out <= 16'h80BF	;
				14'b10111011101000: Data_out <= 16'h80BE	;
				14'b10111011101001: Data_out <= 16'h80BC	;
				14'b10111011101010: Data_out <= 16'h80BB	;
				14'b10111011101011: Data_out <= 16'h80BA	;
				14'b10111011101100: Data_out <= 16'h80B8	;
				14'b10111011101101: Data_out <= 16'h80B7	;
				14'b10111011101110: Data_out <= 16'h80B6	;
				14'b10111011101111: Data_out <= 16'h80B5	;
				14'b10111011110000: Data_out <= 16'h80B3	;
				14'b10111011110001: Data_out <= 16'h80B2	;
				14'b10111011110010: Data_out <= 16'h80B1	;
				14'b10111011110011: Data_out <= 16'h80AF	;
				14'b10111011110100: Data_out <= 16'h80AE	;
				14'b10111011110101: Data_out <= 16'h80AD	;
				14'b10111011110110: Data_out <= 16'h80AB	;
				14'b10111011110111: Data_out <= 16'h80AA	;
				14'b10111011111000: Data_out <= 16'h80A9	;
				14'b10111011111001: Data_out <= 16'h80A8	;
				14'b10111011111010: Data_out <= 16'h80A6	;
				14'b10111011111011: Data_out <= 16'h80A5	;
				14'b10111011111100: Data_out <= 16'h80A4	;
				14'b10111011111101: Data_out <= 16'h80A3	;
				14'b10111011111110: Data_out <= 16'h80A1	;
				14'b10111011111111: Data_out <= 16'h80A0	;
				14'b10111100000000: Data_out <= 16'h809F	;
				14'b10111100000001: Data_out <= 16'h809E	;
				14'b10111100000010: Data_out <= 16'h809C	;
				14'b10111100000011: Data_out <= 16'h809B	;
				14'b10111100000100: Data_out <= 16'h809A	;
				14'b10111100000101: Data_out <= 16'h8099	;
				14'b10111100000110: Data_out <= 16'h8098	;
				14'b10111100000111: Data_out <= 16'h8096	;
				14'b10111100001000: Data_out <= 16'h8095	;
				14'b10111100001001: Data_out <= 16'h8094	;
				14'b10111100001010: Data_out <= 16'h8093	;
				14'b10111100001011: Data_out <= 16'h8092	;
				14'b10111100001100: Data_out <= 16'h8090	;
				14'b10111100001101: Data_out <= 16'h808F	;
				14'b10111100001110: Data_out <= 16'h808E	;
				14'b10111100001111: Data_out <= 16'h808D	;
				14'b10111100010000: Data_out <= 16'h808C	;
				14'b10111100010001: Data_out <= 16'h808B	;
				14'b10111100010010: Data_out <= 16'h8089	;
				14'b10111100010011: Data_out <= 16'h8088	;
				14'b10111100010100: Data_out <= 16'h8087	;
				14'b10111100010101: Data_out <= 16'h8086	;
				14'b10111100010110: Data_out <= 16'h8085	;
				14'b10111100010111: Data_out <= 16'h8084	;
				14'b10111100011000: Data_out <= 16'h8083	;
				14'b10111100011001: Data_out <= 16'h8082	;
				14'b10111100011010: Data_out <= 16'h8080	;
				14'b10111100011011: Data_out <= 16'h807F	;
				14'b10111100011100: Data_out <= 16'h807E	;
				14'b10111100011101: Data_out <= 16'h807D	;
				14'b10111100011110: Data_out <= 16'h807C	;
				14'b10111100011111: Data_out <= 16'h807B	;
				14'b10111100100000: Data_out <= 16'h807A	;
				14'b10111100100001: Data_out <= 16'h8079	;
				14'b10111100100010: Data_out <= 16'h8078	;
				14'b10111100100011: Data_out <= 16'h8077	;
				14'b10111100100100: Data_out <= 16'h8076	;
				14'b10111100100101: Data_out <= 16'h8075	;
				14'b10111100100110: Data_out <= 16'h8074	;
				14'b10111100100111: Data_out <= 16'h8072	;
				14'b10111100101000: Data_out <= 16'h8071	;
				14'b10111100101001: Data_out <= 16'h8070	;
				14'b10111100101010: Data_out <= 16'h806F	;
				14'b10111100101011: Data_out <= 16'h806E	;
				14'b10111100101100: Data_out <= 16'h806D	;
				14'b10111100101101: Data_out <= 16'h806C	;
				14'b10111100101110: Data_out <= 16'h806B	;
				14'b10111100101111: Data_out <= 16'h806A	;
				14'b10111100110000: Data_out <= 16'h8069	;
				14'b10111100110001: Data_out <= 16'h8068	;
				14'b10111100110010: Data_out <= 16'h8067	;
				14'b10111100110011: Data_out <= 16'h8066	;
				14'b10111100110100: Data_out <= 16'h8065	;
				14'b10111100110101: Data_out <= 16'h8064	;
				14'b10111100110110: Data_out <= 16'h8063	;
				14'b10111100110111: Data_out <= 16'h8062	;
				14'b10111100111000: Data_out <= 16'h8061	;
				14'b10111100111001: Data_out <= 16'h8060	;
				14'b10111100111010: Data_out <= 16'h8060	;
				14'b10111100111011: Data_out <= 16'h805F	;
				14'b10111100111100: Data_out <= 16'h805E	;
				14'b10111100111101: Data_out <= 16'h805D	;
				14'b10111100111110: Data_out <= 16'h805C	;
				14'b10111100111111: Data_out <= 16'h805B	;
				14'b10111101000000: Data_out <= 16'h805A	;
				14'b10111101000001: Data_out <= 16'h8059	;
				14'b10111101000010: Data_out <= 16'h8058	;
				14'b10111101000011: Data_out <= 16'h8057	;
				14'b10111101000100: Data_out <= 16'h8056	;
				14'b10111101000101: Data_out <= 16'h8055	;
				14'b10111101000110: Data_out <= 16'h8054	;
				14'b10111101000111: Data_out <= 16'h8054	;
				14'b10111101001000: Data_out <= 16'h8053	;
				14'b10111101001001: Data_out <= 16'h8052	;
				14'b10111101001010: Data_out <= 16'h8051	;
				14'b10111101001011: Data_out <= 16'h8050	;
				14'b10111101001100: Data_out <= 16'h804F	;
				14'b10111101001101: Data_out <= 16'h804E	;
				14'b10111101001110: Data_out <= 16'h804D	;
				14'b10111101001111: Data_out <= 16'h804D	;
				14'b10111101010000: Data_out <= 16'h804C	;
				14'b10111101010001: Data_out <= 16'h804B	;
				14'b10111101010010: Data_out <= 16'h804A	;
				14'b10111101010011: Data_out <= 16'h8049	;
				14'b10111101010100: Data_out <= 16'h8048	;
				14'b10111101010101: Data_out <= 16'h8048	;
				14'b10111101010110: Data_out <= 16'h8047	;
				14'b10111101010111: Data_out <= 16'h8046	;
				14'b10111101011000: Data_out <= 16'h8045	;
				14'b10111101011001: Data_out <= 16'h8044	;
				14'b10111101011010: Data_out <= 16'h8043	;
				14'b10111101011011: Data_out <= 16'h8043	;
				14'b10111101011100: Data_out <= 16'h8042	;
				14'b10111101011101: Data_out <= 16'h8041	;
				14'b10111101011110: Data_out <= 16'h8040	;
				14'b10111101011111: Data_out <= 16'h8040	;
				14'b10111101100000: Data_out <= 16'h803F	;
				14'b10111101100001: Data_out <= 16'h803E	;
				14'b10111101100010: Data_out <= 16'h803D	;
				14'b10111101100011: Data_out <= 16'h803C	;
				14'b10111101100100: Data_out <= 16'h803C	;
				14'b10111101100101: Data_out <= 16'h803B	;
				14'b10111101100110: Data_out <= 16'h803A	;
				14'b10111101100111: Data_out <= 16'h8039	;
				14'b10111101101000: Data_out <= 16'h8039	;
				14'b10111101101001: Data_out <= 16'h8038	;
				14'b10111101101010: Data_out <= 16'h8037	;
				14'b10111101101011: Data_out <= 16'h8037	;
				14'b10111101101100: Data_out <= 16'h8036	;
				14'b10111101101101: Data_out <= 16'h8035	;
				14'b10111101101110: Data_out <= 16'h8034	;
				14'b10111101101111: Data_out <= 16'h8034	;
				14'b10111101110000: Data_out <= 16'h8033	;
				14'b10111101110001: Data_out <= 16'h8032	;
				14'b10111101110010: Data_out <= 16'h8032	;
				14'b10111101110011: Data_out <= 16'h8031	;
				14'b10111101110100: Data_out <= 16'h8030	;
				14'b10111101110101: Data_out <= 16'h8030	;
				14'b10111101110110: Data_out <= 16'h802F	;
				14'b10111101110111: Data_out <= 16'h802E	;
				14'b10111101111000: Data_out <= 16'h802E	;
				14'b10111101111001: Data_out <= 16'h802D	;
				14'b10111101111010: Data_out <= 16'h802C	;
				14'b10111101111011: Data_out <= 16'h802C	;
				14'b10111101111100: Data_out <= 16'h802B	;
				14'b10111101111101: Data_out <= 16'h802A	;
				14'b10111101111110: Data_out <= 16'h802A	;
				14'b10111101111111: Data_out <= 16'h8029	;
				14'b10111110000000: Data_out <= 16'h8029	;
				14'b10111110000001: Data_out <= 16'h8028	;
				14'b10111110000010: Data_out <= 16'h8027	;
				14'b10111110000011: Data_out <= 16'h8027	;
				14'b10111110000100: Data_out <= 16'h8026	;
				14'b10111110000101: Data_out <= 16'h8026	;
				14'b10111110000110: Data_out <= 16'h8025	;
				14'b10111110000111: Data_out <= 16'h8024	;
				14'b10111110001000: Data_out <= 16'h8024	;
				14'b10111110001001: Data_out <= 16'h8023	;
				14'b10111110001010: Data_out <= 16'h8023	;
				14'b10111110001011: Data_out <= 16'h8022	;
				14'b10111110001100: Data_out <= 16'h8022	;
				14'b10111110001101: Data_out <= 16'h8021	;
				14'b10111110001110: Data_out <= 16'h8020	;
				14'b10111110001111: Data_out <= 16'h8020	;
				14'b10111110010000: Data_out <= 16'h801F	;
				14'b10111110010001: Data_out <= 16'h801F	;
				14'b10111110010010: Data_out <= 16'h801E	;
				14'b10111110010011: Data_out <= 16'h801E	;
				14'b10111110010100: Data_out <= 16'h801D	;
				14'b10111110010101: Data_out <= 16'h801D	;
				14'b10111110010110: Data_out <= 16'h801C	;
				14'b10111110010111: Data_out <= 16'h801C	;
				14'b10111110011000: Data_out <= 16'h801B	;
				14'b10111110011001: Data_out <= 16'h801B	;
				14'b10111110011010: Data_out <= 16'h801A	;
				14'b10111110011011: Data_out <= 16'h801A	;
				14'b10111110011100: Data_out <= 16'h8019	;
				14'b10111110011101: Data_out <= 16'h8019	;
				14'b10111110011110: Data_out <= 16'h8018	;
				14'b10111110011111: Data_out <= 16'h8018	;
				14'b10111110100000: Data_out <= 16'h8017	;
				14'b10111110100001: Data_out <= 16'h8017	;
				14'b10111110100010: Data_out <= 16'h8016	;
				14'b10111110100011: Data_out <= 16'h8016	;
				14'b10111110100100: Data_out <= 16'h8015	;
				14'b10111110100101: Data_out <= 16'h8015	;
				14'b10111110100110: Data_out <= 16'h8015	;
				14'b10111110100111: Data_out <= 16'h8014	;
				14'b10111110101000: Data_out <= 16'h8014	;
				14'b10111110101001: Data_out <= 16'h8013	;
				14'b10111110101010: Data_out <= 16'h8013	;
				14'b10111110101011: Data_out <= 16'h8013	;
				14'b10111110101100: Data_out <= 16'h8012	;
				14'b10111110101101: Data_out <= 16'h8012	;
				14'b10111110101110: Data_out <= 16'h8011	;
				14'b10111110101111: Data_out <= 16'h8011	;
				14'b10111110110000: Data_out <= 16'h8011	;
				14'b10111110110001: Data_out <= 16'h8010	;
				14'b10111110110010: Data_out <= 16'h8010	;
				14'b10111110110011: Data_out <= 16'h800F	;
				14'b10111110110100: Data_out <= 16'h800F	;
				14'b10111110110101: Data_out <= 16'h800F	;
				14'b10111110110110: Data_out <= 16'h800E	;
				14'b10111110110111: Data_out <= 16'h800E	;
				14'b10111110111000: Data_out <= 16'h800E	;
				14'b10111110111001: Data_out <= 16'h800D	;
				14'b10111110111010: Data_out <= 16'h800D	;
				14'b10111110111011: Data_out <= 16'h800D	;
				14'b10111110111100: Data_out <= 16'h800C	;
				14'b10111110111101: Data_out <= 16'h800C	;
				14'b10111110111110: Data_out <= 16'h800C	;
				14'b10111110111111: Data_out <= 16'h800B	;
				14'b10111111000000: Data_out <= 16'h800B	;
				14'b10111111000001: Data_out <= 16'h800B	;
				14'b10111111000010: Data_out <= 16'h800A	;
				14'b10111111000011: Data_out <= 16'h800A	;
				14'b10111111000100: Data_out <= 16'h800A	;
				14'b10111111000101: Data_out <= 16'h8009	;
				14'b10111111000110: Data_out <= 16'h8009	;
				14'b10111111000111: Data_out <= 16'h8009	;
				14'b10111111001000: Data_out <= 16'h8009	;
				14'b10111111001001: Data_out <= 16'h8008	;
				14'b10111111001010: Data_out <= 16'h8008	;
				14'b10111111001011: Data_out <= 16'h8008	;
				14'b10111111001100: Data_out <= 16'h8008	;
				14'b10111111001101: Data_out <= 16'h8007	;
				14'b10111111001110: Data_out <= 16'h8007	;
				14'b10111111001111: Data_out <= 16'h8007	;
				14'b10111111010000: Data_out <= 16'h8007	;
				14'b10111111010001: Data_out <= 16'h8006	;
				14'b10111111010010: Data_out <= 16'h8006	;
				14'b10111111010011: Data_out <= 16'h8006	;
				14'b10111111010100: Data_out <= 16'h8006	;
				14'b10111111010101: Data_out <= 16'h8006	;
				14'b10111111010110: Data_out <= 16'h8005	;
				14'b10111111010111: Data_out <= 16'h8005	;
				14'b10111111011000: Data_out <= 16'h8005	;
				14'b10111111011001: Data_out <= 16'h8005	;
				14'b10111111011010: Data_out <= 16'h8005	;
				14'b10111111011011: Data_out <= 16'h8004	;
				14'b10111111011100: Data_out <= 16'h8004	;
				14'b10111111011101: Data_out <= 16'h8004	;
				14'b10111111011110: Data_out <= 16'h8004	;
				14'b10111111011111: Data_out <= 16'h8004	;
				14'b10111111100000: Data_out <= 16'h8004	;
				14'b10111111100001: Data_out <= 16'h8003	;
				14'b10111111100010: Data_out <= 16'h8003	;
				14'b10111111100011: Data_out <= 16'h8003	;
				14'b10111111100100: Data_out <= 16'h8003	;
				14'b10111111100101: Data_out <= 16'h8003	;
				14'b10111111100110: Data_out <= 16'h8003	;
				14'b10111111100111: Data_out <= 16'h8003	;
				14'b10111111101000: Data_out <= 16'h8002	;
				14'b10111111101001: Data_out <= 16'h8002	;
				14'b10111111101010: Data_out <= 16'h8002	;
				14'b10111111101011: Data_out <= 16'h8002	;
				14'b10111111101100: Data_out <= 16'h8002	;
				14'b10111111101101: Data_out <= 16'h8002	;
				14'b10111111101110: Data_out <= 16'h8002	;
				14'b10111111101111: Data_out <= 16'h8002	;
				14'b10111111110000: Data_out <= 16'h8002	;
				14'b10111111110001: Data_out <= 16'h8002	;
				14'b10111111110010: Data_out <= 16'h8002	;
				14'b10111111110011: Data_out <= 16'h8002	;
				14'b10111111110100: Data_out <= 16'h8001	;
				14'b10111111110101: Data_out <= 16'h8001	;
				14'b10111111110110: Data_out <= 16'h8001	;
				14'b10111111110111: Data_out <= 16'h8001	;
				14'b10111111111000: Data_out <= 16'h8001	;
				14'b10111111111001: Data_out <= 16'h8001	;
				14'b10111111111010: Data_out <= 16'h8001	;
				14'b10111111111011: Data_out <= 16'h8001	;
				14'b10111111111100: Data_out <= 16'h8001	;
				14'b10111111111101: Data_out <= 16'h8001	;
				14'b10111111111110: Data_out <= 16'h8001	;
				14'b10111111111111: Data_out <= 16'h8001	;
				/////////////////////////////////////////////////////////////////////////////////////////////
				//	negative	half-cycle of rise......
				14'b11000000000000: Data_out <= 16'h8001	;
				14'b11000000000001: Data_out <= 16'h8001	;
				14'b11000000000010: Data_out <= 16'h8001	;
				14'b11000000000011: Data_out <= 16'h8001	;
				14'b11000000000100: Data_out <= 16'h8001	;
				14'b11000000000101: Data_out <= 16'h8001	;
				14'b11000000000110: Data_out <= 16'h8001	;
				14'b11000000000111: Data_out <= 16'h8001	;
				14'b11000000001000: Data_out <= 16'h8001	;
				14'b11000000001001: Data_out <= 16'h8001	;
				14'b11000000001010: Data_out <= 16'h8001	;
				14'b11000000001011: Data_out <= 16'h8001	;
				14'b11000000001100: Data_out <= 16'h8001	;
				14'b11000000001101: Data_out <= 16'h8002	;
				14'b11000000001110: Data_out <= 16'h8002	;
				14'b11000000001111: Data_out <= 16'h8002	;
				14'b11000000010000: Data_out <= 16'h8002	;
				14'b11000000010001: Data_out <= 16'h8002	;
				14'b11000000010010: Data_out <= 16'h8002	;
				14'b11000000010011: Data_out <= 16'h8002	;
				14'b11000000010100: Data_out <= 16'h8002	;
				14'b11000000010101: Data_out <= 16'h8002	;
				14'b11000000010110: Data_out <= 16'h8002	;
				14'b11000000010111: Data_out <= 16'h8002	;
				14'b11000000011000: Data_out <= 16'h8002	;
				14'b11000000011001: Data_out <= 16'h8003	;
				14'b11000000011010: Data_out <= 16'h8003	;
				14'b11000000011011: Data_out <= 16'h8003	;
				14'b11000000011100: Data_out <= 16'h8003	;
				14'b11000000011101: Data_out <= 16'h8003	;
				14'b11000000011110: Data_out <= 16'h8003	;
				14'b11000000011111: Data_out <= 16'h8003	;
				14'b11000000100000: Data_out <= 16'h8004	;
				14'b11000000100001: Data_out <= 16'h8004	;
				14'b11000000100010: Data_out <= 16'h8004	;
				14'b11000000100011: Data_out <= 16'h8004	;
				14'b11000000100100: Data_out <= 16'h8004	;
				14'b11000000100101: Data_out <= 16'h8004	;
				14'b11000000100110: Data_out <= 16'h8005	;
				14'b11000000100111: Data_out <= 16'h8005	;
				14'b11000000101000: Data_out <= 16'h8005	;
				14'b11000000101001: Data_out <= 16'h8005	;
				14'b11000000101010: Data_out <= 16'h8005	;
				14'b11000000101011: Data_out <= 16'h8006	;
				14'b11000000101100: Data_out <= 16'h8006	;
				14'b11000000101101: Data_out <= 16'h8006	;
				14'b11000000101110: Data_out <= 16'h8006	;
				14'b11000000101111: Data_out <= 16'h8006	;
				14'b11000000110000: Data_out <= 16'h8007	;
				14'b11000000110001: Data_out <= 16'h8007	;
				14'b11000000110010: Data_out <= 16'h8007	;
				14'b11000000110011: Data_out <= 16'h8007	;
				14'b11000000110100: Data_out <= 16'h8008	;
				14'b11000000110101: Data_out <= 16'h8008	;
				14'b11000000110110: Data_out <= 16'h8008	;
				14'b11000000110111: Data_out <= 16'h8008	;
				14'b11000000111000: Data_out <= 16'h8009	;
				14'b11000000111001: Data_out <= 16'h8009	;
				14'b11000000111010: Data_out <= 16'h8009	;
				14'b11000000111011: Data_out <= 16'h8009	;
				14'b11000000111100: Data_out <= 16'h800A	;
				14'b11000000111101: Data_out <= 16'h800A	;
				14'b11000000111110: Data_out <= 16'h800A	;
				14'b11000000111111: Data_out <= 16'h800B	;
				14'b11000001000000: Data_out <= 16'h800B	;
				14'b11000001000001: Data_out <= 16'h800B	;
				14'b11000001000010: Data_out <= 16'h800C	;
				14'b11000001000011: Data_out <= 16'h800C	;
				14'b11000001000100: Data_out <= 16'h800C	;
				14'b11000001000101: Data_out <= 16'h800D	;
				14'b11000001000110: Data_out <= 16'h800D	;
				14'b11000001000111: Data_out <= 16'h800D	;
				14'b11000001001000: Data_out <= 16'h800E	;
				14'b11000001001001: Data_out <= 16'h800E	;
				14'b11000001001010: Data_out <= 16'h800E	;
				14'b11000001001011: Data_out <= 16'h800F	;
				14'b11000001001100: Data_out <= 16'h800F	;
				14'b11000001001101: Data_out <= 16'h800F	;
				14'b11000001001110: Data_out <= 16'h8010	;
				14'b11000001001111: Data_out <= 16'h8010	;
				14'b11000001010000: Data_out <= 16'h8011	;
				14'b11000001010001: Data_out <= 16'h8011	;
				14'b11000001010010: Data_out <= 16'h8011	;
				14'b11000001010011: Data_out <= 16'h8012	;
				14'b11000001010100: Data_out <= 16'h8012	;
				14'b11000001010101: Data_out <= 16'h8013	;
				14'b11000001010110: Data_out <= 16'h8013	;
				14'b11000001010111: Data_out <= 16'h8013	;
				14'b11000001011000: Data_out <= 16'h8014	;
				14'b11000001011001: Data_out <= 16'h8014	;
				14'b11000001011010: Data_out <= 16'h8015	;
				14'b11000001011011: Data_out <= 16'h8015	;
				14'b11000001011100: Data_out <= 16'h8015	;
				14'b11000001011101: Data_out <= 16'h8016	;
				14'b11000001011110: Data_out <= 16'h8016	;
				14'b11000001011111: Data_out <= 16'h8017	;
				14'b11000001100000: Data_out <= 16'h8017	;
				14'b11000001100001: Data_out <= 16'h8018	;
				14'b11000001100010: Data_out <= 16'h8018	;
				14'b11000001100011: Data_out <= 16'h8019	;
				14'b11000001100100: Data_out <= 16'h8019	;
				14'b11000001100101: Data_out <= 16'h801A	;
				14'b11000001100110: Data_out <= 16'h801A	;
				14'b11000001100111: Data_out <= 16'h801B	;
				14'b11000001101000: Data_out <= 16'h801B	;
				14'b11000001101001: Data_out <= 16'h801C	;
				14'b11000001101010: Data_out <= 16'h801C	;
				14'b11000001101011: Data_out <= 16'h801D	;
				14'b11000001101100: Data_out <= 16'h801D	;
				14'b11000001101101: Data_out <= 16'h801E	;
				14'b11000001101110: Data_out <= 16'h801E	;
				14'b11000001101111: Data_out <= 16'h801F	;
				14'b11000001110000: Data_out <= 16'h801F	;
				14'b11000001110001: Data_out <= 16'h8020	;
				14'b11000001110010: Data_out <= 16'h8020	;
				14'b11000001110011: Data_out <= 16'h8021	;
				14'b11000001110100: Data_out <= 16'h8022	;
				14'b11000001110101: Data_out <= 16'h8022	;
				14'b11000001110110: Data_out <= 16'h8023	;
				14'b11000001110111: Data_out <= 16'h8023	;
				14'b11000001111000: Data_out <= 16'h8024	;
				14'b11000001111001: Data_out <= 16'h8024	;
				14'b11000001111010: Data_out <= 16'h8025	;
				14'b11000001111011: Data_out <= 16'h8026	;
				14'b11000001111100: Data_out <= 16'h8026	;
				14'b11000001111101: Data_out <= 16'h8027	;
				14'b11000001111110: Data_out <= 16'h8027	;
				14'b11000001111111: Data_out <= 16'h8028	;
				14'b11000010000000: Data_out <= 16'h8029	;
				14'b11000010000001: Data_out <= 16'h8029	;
				14'b11000010000010: Data_out <= 16'h802A	;
				14'b11000010000011: Data_out <= 16'h802A	;
				14'b11000010000100: Data_out <= 16'h802B	;
				14'b11000010000101: Data_out <= 16'h802C	;
				14'b11000010000110: Data_out <= 16'h802C	;
				14'b11000010000111: Data_out <= 16'h802D	;
				14'b11000010001000: Data_out <= 16'h802E	;
				14'b11000010001001: Data_out <= 16'h802E	;
				14'b11000010001010: Data_out <= 16'h802F	;
				14'b11000010001011: Data_out <= 16'h8030	;
				14'b11000010001100: Data_out <= 16'h8030	;
				14'b11000010001101: Data_out <= 16'h8031	;
				14'b11000010001110: Data_out <= 16'h8032	;
				14'b11000010001111: Data_out <= 16'h8032	;
				14'b11000010010000: Data_out <= 16'h8033	;
				14'b11000010010001: Data_out <= 16'h8034	;
				14'b11000010010010: Data_out <= 16'h8034	;
				14'b11000010010011: Data_out <= 16'h8035	;
				14'b11000010010100: Data_out <= 16'h8036	;
				14'b11000010010101: Data_out <= 16'h8037	;
				14'b11000010010110: Data_out <= 16'h8037	;
				14'b11000010010111: Data_out <= 16'h8038	;
				14'b11000010011000: Data_out <= 16'h8039	;
				14'b11000010011001: Data_out <= 16'h8039	;
				14'b11000010011010: Data_out <= 16'h803A	;
				14'b11000010011011: Data_out <= 16'h803B	;
				14'b11000010011100: Data_out <= 16'h803C	;
				14'b11000010011101: Data_out <= 16'h803C	;
				14'b11000010011110: Data_out <= 16'h803D	;
				14'b11000010011111: Data_out <= 16'h803E	;
				14'b11000010100000: Data_out <= 16'h803F	;
				14'b11000010100001: Data_out <= 16'h8040	;
				14'b11000010100010: Data_out <= 16'h8040	;
				14'b11000010100011: Data_out <= 16'h8041	;
				14'b11000010100100: Data_out <= 16'h8042	;
				14'b11000010100101: Data_out <= 16'h8043	;
				14'b11000010100110: Data_out <= 16'h8043	;
				14'b11000010100111: Data_out <= 16'h8044	;
				14'b11000010101000: Data_out <= 16'h8045	;
				14'b11000010101001: Data_out <= 16'h8046	;
				14'b11000010101010: Data_out <= 16'h8047	;
				14'b11000010101011: Data_out <= 16'h8048	;
				14'b11000010101100: Data_out <= 16'h8048	;
				14'b11000010101101: Data_out <= 16'h8049	;
				14'b11000010101110: Data_out <= 16'h804A	;
				14'b11000010101111: Data_out <= 16'h804B	;
				14'b11000010110000: Data_out <= 16'h804C	;
				14'b11000010110001: Data_out <= 16'h804D	;
				14'b11000010110010: Data_out <= 16'h804D	;
				14'b11000010110011: Data_out <= 16'h804E	;
				14'b11000010110100: Data_out <= 16'h804F	;
				14'b11000010110101: Data_out <= 16'h8050	;
				14'b11000010110110: Data_out <= 16'h8051	;
				14'b11000010110111: Data_out <= 16'h8052	;
				14'b11000010111000: Data_out <= 16'h8053	;
				14'b11000010111001: Data_out <= 16'h8054	;
				14'b11000010111010: Data_out <= 16'h8054	;
				14'b11000010111011: Data_out <= 16'h8055	;
				14'b11000010111100: Data_out <= 16'h8056	;
				14'b11000010111101: Data_out <= 16'h8057	;
				14'b11000010111110: Data_out <= 16'h8058	;
				14'b11000010111111: Data_out <= 16'h8059	;
				14'b11000011000000: Data_out <= 16'h805A	;
				14'b11000011000001: Data_out <= 16'h805B	;
				14'b11000011000010: Data_out <= 16'h805C	;
				14'b11000011000011: Data_out <= 16'h805D	;
				14'b11000011000100: Data_out <= 16'h805E	;
				14'b11000011000101: Data_out <= 16'h805F	;
				14'b11000011000110: Data_out <= 16'h8060	;
				14'b11000011000111: Data_out <= 16'h8060	;
				14'b11000011001000: Data_out <= 16'h8061	;
				14'b11000011001001: Data_out <= 16'h8062	;
				14'b11000011001010: Data_out <= 16'h8063	;
				14'b11000011001011: Data_out <= 16'h8064	;
				14'b11000011001100: Data_out <= 16'h8065	;
				14'b11000011001101: Data_out <= 16'h8066	;
				14'b11000011001110: Data_out <= 16'h8067	;
				14'b11000011001111: Data_out <= 16'h8068	;
				14'b11000011010000: Data_out <= 16'h8069	;
				14'b11000011010001: Data_out <= 16'h806A	;
				14'b11000011010010: Data_out <= 16'h806B	;
				14'b11000011010011: Data_out <= 16'h806C	;
				14'b11000011010100: Data_out <= 16'h806D	;
				14'b11000011010101: Data_out <= 16'h806E	;
				14'b11000011010110: Data_out <= 16'h806F	;
				14'b11000011010111: Data_out <= 16'h8070	;
				14'b11000011011000: Data_out <= 16'h8071	;
				14'b11000011011001: Data_out <= 16'h8072	;
				14'b11000011011010: Data_out <= 16'h8074	;
				14'b11000011011011: Data_out <= 16'h8075	;
				14'b11000011011100: Data_out <= 16'h8076	;
				14'b11000011011101: Data_out <= 16'h8077	;
				14'b11000011011110: Data_out <= 16'h8078	;
				14'b11000011011111: Data_out <= 16'h8079	;
				14'b11000011100000: Data_out <= 16'h807A	;
				14'b11000011100001: Data_out <= 16'h807B	;
				14'b11000011100010: Data_out <= 16'h807C	;
				14'b11000011100011: Data_out <= 16'h807D	;
				14'b11000011100100: Data_out <= 16'h807E	;
				14'b11000011100101: Data_out <= 16'h807F	;
				14'b11000011100110: Data_out <= 16'h8080	;
				14'b11000011100111: Data_out <= 16'h8082	;
				14'b11000011101000: Data_out <= 16'h8083	;
				14'b11000011101001: Data_out <= 16'h8084	;
				14'b11000011101010: Data_out <= 16'h8085	;
				14'b11000011101011: Data_out <= 16'h8086	;
				14'b11000011101100: Data_out <= 16'h8087	;
				14'b11000011101101: Data_out <= 16'h8088	;
				14'b11000011101110: Data_out <= 16'h8089	;
				14'b11000011101111: Data_out <= 16'h808B	;
				14'b11000011110000: Data_out <= 16'h808C	;
				14'b11000011110001: Data_out <= 16'h808D	;
				14'b11000011110010: Data_out <= 16'h808E	;
				14'b11000011110011: Data_out <= 16'h808F	;
				14'b11000011110100: Data_out <= 16'h8090	;
				14'b11000011110101: Data_out <= 16'h8092	;
				14'b11000011110110: Data_out <= 16'h8093	;
				14'b11000011110111: Data_out <= 16'h8094	;
				14'b11000011111000: Data_out <= 16'h8095	;
				14'b11000011111001: Data_out <= 16'h8096	;
				14'b11000011111010: Data_out <= 16'h8098	;
				14'b11000011111011: Data_out <= 16'h8099	;
				14'b11000011111100: Data_out <= 16'h809A	;
				14'b11000011111101: Data_out <= 16'h809B	;
				14'b11000011111110: Data_out <= 16'h809C	;
				14'b11000011111111: Data_out <= 16'h809E	;
				14'b11000100000000: Data_out <= 16'h809F	;
				14'b11000100000001: Data_out <= 16'h80A0	;
				14'b11000100000010: Data_out <= 16'h80A1	;
				14'b11000100000011: Data_out <= 16'h80A3	;
				14'b11000100000100: Data_out <= 16'h80A4	;
				14'b11000100000101: Data_out <= 16'h80A5	;
				14'b11000100000110: Data_out <= 16'h80A6	;
				14'b11000100000111: Data_out <= 16'h80A8	;
				14'b11000100001000: Data_out <= 16'h80A9	;
				14'b11000100001001: Data_out <= 16'h80AA	;
				14'b11000100001010: Data_out <= 16'h80AB	;
				14'b11000100001011: Data_out <= 16'h80AD	;
				14'b11000100001100: Data_out <= 16'h80AE	;
				14'b11000100001101: Data_out <= 16'h80AF	;
				14'b11000100001110: Data_out <= 16'h80B1	;
				14'b11000100001111: Data_out <= 16'h80B2	;
				14'b11000100010000: Data_out <= 16'h80B3	;
				14'b11000100010001: Data_out <= 16'h80B5	;
				14'b11000100010010: Data_out <= 16'h80B6	;
				14'b11000100010011: Data_out <= 16'h80B7	;
				14'b11000100010100: Data_out <= 16'h80B8	;
				14'b11000100010101: Data_out <= 16'h80BA	;
				14'b11000100010110: Data_out <= 16'h80BB	;
				14'b11000100010111: Data_out <= 16'h80BC	;
				14'b11000100011000: Data_out <= 16'h80BE	;
				14'b11000100011001: Data_out <= 16'h80BF	;
				14'b11000100011010: Data_out <= 16'h80C1	;
				14'b11000100011011: Data_out <= 16'h80C2	;
				14'b11000100011100: Data_out <= 16'h80C3	;
				14'b11000100011101: Data_out <= 16'h80C5	;
				14'b11000100011110: Data_out <= 16'h80C6	;
				14'b11000100011111: Data_out <= 16'h80C7	;
				14'b11000100100000: Data_out <= 16'h80C9	;
				14'b11000100100001: Data_out <= 16'h80CA	;
				14'b11000100100010: Data_out <= 16'h80CC	;
				14'b11000100100011: Data_out <= 16'h80CD	;
				14'b11000100100100: Data_out <= 16'h80CE	;
				14'b11000100100101: Data_out <= 16'h80D0	;
				14'b11000100100110: Data_out <= 16'h80D1	;
				14'b11000100100111: Data_out <= 16'h80D3	;
				14'b11000100101000: Data_out <= 16'h80D4	;
				14'b11000100101001: Data_out <= 16'h80D5	;
				14'b11000100101010: Data_out <= 16'h80D7	;
				14'b11000100101011: Data_out <= 16'h80D8	;
				14'b11000100101100: Data_out <= 16'h80DA	;
				14'b11000100101101: Data_out <= 16'h80DB	;
				14'b11000100101110: Data_out <= 16'h80DD	;
				14'b11000100101111: Data_out <= 16'h80DE	;
				14'b11000100110000: Data_out <= 16'h80E0	;
				14'b11000100110001: Data_out <= 16'h80E1	;
				14'b11000100110010: Data_out <= 16'h80E2	;
				14'b11000100110011: Data_out <= 16'h80E4	;
				14'b11000100110100: Data_out <= 16'h80E5	;
				14'b11000100110101: Data_out <= 16'h80E7	;
				14'b11000100110110: Data_out <= 16'h80E8	;
				14'b11000100110111: Data_out <= 16'h80EA	;
				14'b11000100111000: Data_out <= 16'h80EB	;
				14'b11000100111001: Data_out <= 16'h80ED	;
				14'b11000100111010: Data_out <= 16'h80EE	;
				14'b11000100111011: Data_out <= 16'h80F0	;
				14'b11000100111100: Data_out <= 16'h80F1	;
				14'b11000100111101: Data_out <= 16'h80F3	;
				14'b11000100111110: Data_out <= 16'h80F4	;
				14'b11000100111111: Data_out <= 16'h80F6	;
				14'b11000101000000: Data_out <= 16'h80F8	;
				14'b11000101000001: Data_out <= 16'h80F9	;
				14'b11000101000010: Data_out <= 16'h80FB	;
				14'b11000101000011: Data_out <= 16'h80FC	;
				14'b11000101000100: Data_out <= 16'h80FE	;
				14'b11000101000101: Data_out <= 16'h80FF	;
				14'b11000101000110: Data_out <= 16'h8101	;
				14'b11000101000111: Data_out <= 16'h8102	;
				14'b11000101001000: Data_out <= 16'h8104	;
				14'b11000101001001: Data_out <= 16'h8106	;
				14'b11000101001010: Data_out <= 16'h8107	;
				14'b11000101001011: Data_out <= 16'h8109	;
				14'b11000101001100: Data_out <= 16'h810A	;
				14'b11000101001101: Data_out <= 16'h810C	;
				14'b11000101001110: Data_out <= 16'h810E	;
				14'b11000101001111: Data_out <= 16'h810F	;
				14'b11000101010000: Data_out <= 16'h8111	;
				14'b11000101010001: Data_out <= 16'h8112	;
				14'b11000101010010: Data_out <= 16'h8114	;
				14'b11000101010011: Data_out <= 16'h8116	;
				14'b11000101010100: Data_out <= 16'h8117	;
				14'b11000101010101: Data_out <= 16'h8119	;
				14'b11000101010110: Data_out <= 16'h811B	;
				14'b11000101010111: Data_out <= 16'h811C	;
				14'b11000101011000: Data_out <= 16'h811E	;
				14'b11000101011001: Data_out <= 16'h811F	;
				14'b11000101011010: Data_out <= 16'h8121	;
				14'b11000101011011: Data_out <= 16'h8123	;
				14'b11000101011100: Data_out <= 16'h8124	;
				14'b11000101011101: Data_out <= 16'h8126	;
				14'b11000101011110: Data_out <= 16'h8128	;
				14'b11000101011111: Data_out <= 16'h812A	;
				14'b11000101100000: Data_out <= 16'h812B	;
				14'b11000101100001: Data_out <= 16'h812D	;
				14'b11000101100010: Data_out <= 16'h812F	;
				14'b11000101100011: Data_out <= 16'h8130	;
				14'b11000101100100: Data_out <= 16'h8132	;
				14'b11000101100101: Data_out <= 16'h8134	;
				14'b11000101100110: Data_out <= 16'h8135	;
				14'b11000101100111: Data_out <= 16'h8137	;
				14'b11000101101000: Data_out <= 16'h8139	;
				14'b11000101101001: Data_out <= 16'h813B	;
				14'b11000101101010: Data_out <= 16'h813C	;
				14'b11000101101011: Data_out <= 16'h813E	;
				14'b11000101101100: Data_out <= 16'h8140	;
				14'b11000101101101: Data_out <= 16'h8142	;
				14'b11000101101110: Data_out <= 16'h8143	;
				14'b11000101101111: Data_out <= 16'h8145	;
				14'b11000101110000: Data_out <= 16'h8147	;
				14'b11000101110001: Data_out <= 16'h8149	;
				14'b11000101110010: Data_out <= 16'h814A	;
				14'b11000101110011: Data_out <= 16'h814C	;
				14'b11000101110100: Data_out <= 16'h814E	;
				14'b11000101110101: Data_out <= 16'h8150	;
				14'b11000101110110: Data_out <= 16'h8152	;
				14'b11000101110111: Data_out <= 16'h8153	;
				14'b11000101111000: Data_out <= 16'h8155	;
				14'b11000101111001: Data_out <= 16'h8157	;
				14'b11000101111010: Data_out <= 16'h8159	;
				14'b11000101111011: Data_out <= 16'h815B	;
				14'b11000101111100: Data_out <= 16'h815C	;
				14'b11000101111101: Data_out <= 16'h815E	;
				14'b11000101111110: Data_out <= 16'h8160	;
				14'b11000101111111: Data_out <= 16'h8162	;
				14'b11000110000000: Data_out <= 16'h8164	;
				14'b11000110000001: Data_out <= 16'h8166	;
				14'b11000110000010: Data_out <= 16'h8167	;
				14'b11000110000011: Data_out <= 16'h8169	;
				14'b11000110000100: Data_out <= 16'h816B	;
				14'b11000110000101: Data_out <= 16'h816D	;
				14'b11000110000110: Data_out <= 16'h816F	;
				14'b11000110000111: Data_out <= 16'h8171	;
				14'b11000110001000: Data_out <= 16'h8173	;
				14'b11000110001001: Data_out <= 16'h8175	;
				14'b11000110001010: Data_out <= 16'h8176	;
				14'b11000110001011: Data_out <= 16'h8178	;
				14'b11000110001100: Data_out <= 16'h817A	;
				14'b11000110001101: Data_out <= 16'h817C	;
				14'b11000110001110: Data_out <= 16'h817E	;
				14'b11000110001111: Data_out <= 16'h8180	;
				14'b11000110010000: Data_out <= 16'h8182	;
				14'b11000110010001: Data_out <= 16'h8184	;
				14'b11000110010010: Data_out <= 16'h8186	;
				14'b11000110010011: Data_out <= 16'h8188	;
				14'b11000110010100: Data_out <= 16'h818A	;
				14'b11000110010101: Data_out <= 16'h818C	;
				14'b11000110010110: Data_out <= 16'h818D	;
				14'b11000110010111: Data_out <= 16'h818F	;
				14'b11000110011000: Data_out <= 16'h8191	;
				14'b11000110011001: Data_out <= 16'h8193	;
				14'b11000110011010: Data_out <= 16'h8195	;
				14'b11000110011011: Data_out <= 16'h8197	;
				14'b11000110011100: Data_out <= 16'h8199	;
				14'b11000110011101: Data_out <= 16'h819B	;
				14'b11000110011110: Data_out <= 16'h819D	;
				14'b11000110011111: Data_out <= 16'h819F	;
				14'b11000110100000: Data_out <= 16'h81A1	;
				14'b11000110100001: Data_out <= 16'h81A3	;
				14'b11000110100010: Data_out <= 16'h81A5	;
				14'b11000110100011: Data_out <= 16'h81A7	;
				14'b11000110100100: Data_out <= 16'h81A9	;
				14'b11000110100101: Data_out <= 16'h81AB	;
				14'b11000110100110: Data_out <= 16'h81AD	;
				14'b11000110100111: Data_out <= 16'h81AF	;
				14'b11000110101000: Data_out <= 16'h81B1	;
				14'b11000110101001: Data_out <= 16'h81B3	;
				14'b11000110101010: Data_out <= 16'h81B5	;
				14'b11000110101011: Data_out <= 16'h81B7	;
				14'b11000110101100: Data_out <= 16'h81B9	;
				14'b11000110101101: Data_out <= 16'h81BC	;
				14'b11000110101110: Data_out <= 16'h81BE	;
				14'b11000110101111: Data_out <= 16'h81C0	;
				14'b11000110110000: Data_out <= 16'h81C2	;
				14'b11000110110001: Data_out <= 16'h81C4	;
				14'b11000110110010: Data_out <= 16'h81C6	;
				14'b11000110110011: Data_out <= 16'h81C8	;
				14'b11000110110100: Data_out <= 16'h81CA	;
				14'b11000110110101: Data_out <= 16'h81CC	;
				14'b11000110110110: Data_out <= 16'h81CE	;
				14'b11000110110111: Data_out <= 16'h81D0	;
				14'b11000110111000: Data_out <= 16'h81D2	;
				14'b11000110111001: Data_out <= 16'h81D5	;
				14'b11000110111010: Data_out <= 16'h81D7	;
				14'b11000110111011: Data_out <= 16'h81D9	;
				14'b11000110111100: Data_out <= 16'h81DB	;
				14'b11000110111101: Data_out <= 16'h81DD	;
				14'b11000110111110: Data_out <= 16'h81DF	;
				14'b11000110111111: Data_out <= 16'h81E1	;
				14'b11000111000000: Data_out <= 16'h81E4	;
				14'b11000111000001: Data_out <= 16'h81E6	;
				14'b11000111000010: Data_out <= 16'h81E8	;
				14'b11000111000011: Data_out <= 16'h81EA	;
				14'b11000111000100: Data_out <= 16'h81EC	;
				14'b11000111000101: Data_out <= 16'h81EE	;
				14'b11000111000110: Data_out <= 16'h81F0	;
				14'b11000111000111: Data_out <= 16'h81F3	;
				14'b11000111001000: Data_out <= 16'h81F5	;
				14'b11000111001001: Data_out <= 16'h81F7	;
				14'b11000111001010: Data_out <= 16'h81F9	;
				14'b11000111001011: Data_out <= 16'h81FB	;
				14'b11000111001100: Data_out <= 16'h81FE	;
				14'b11000111001101: Data_out <= 16'h8200	;
				14'b11000111001110: Data_out <= 16'h8202	;
				14'b11000111001111: Data_out <= 16'h8204	;
				14'b11000111010000: Data_out <= 16'h8206	;
				14'b11000111010001: Data_out <= 16'h8209	;
				14'b11000111010010: Data_out <= 16'h820B	;
				14'b11000111010011: Data_out <= 16'h820D	;
				14'b11000111010100: Data_out <= 16'h820F	;
				14'b11000111010101: Data_out <= 16'h8212	;
				14'b11000111010110: Data_out <= 16'h8214	;
				14'b11000111010111: Data_out <= 16'h8216	;
				14'b11000111011000: Data_out <= 16'h8218	;
				14'b11000111011001: Data_out <= 16'h821B	;
				14'b11000111011010: Data_out <= 16'h821D	;
				14'b11000111011011: Data_out <= 16'h821F	;
				14'b11000111011100: Data_out <= 16'h8222	;
				14'b11000111011101: Data_out <= 16'h8224	;
				14'b11000111011110: Data_out <= 16'h8226	;
				14'b11000111011111: Data_out <= 16'h8228	;
				14'b11000111100000: Data_out <= 16'h822B	;
				14'b11000111100001: Data_out <= 16'h822D	;
				14'b11000111100010: Data_out <= 16'h822F	;
				14'b11000111100011: Data_out <= 16'h8232	;
				14'b11000111100100: Data_out <= 16'h8234	;
				14'b11000111100101: Data_out <= 16'h8236	;
				14'b11000111100110: Data_out <= 16'h8239	;
				14'b11000111100111: Data_out <= 16'h823B	;
				14'b11000111101000: Data_out <= 16'h823D	;
				14'b11000111101001: Data_out <= 16'h8240	;
				14'b11000111101010: Data_out <= 16'h8242	;
				14'b11000111101011: Data_out <= 16'h8244	;
				14'b11000111101100: Data_out <= 16'h8247	;
				14'b11000111101101: Data_out <= 16'h8249	;
				14'b11000111101110: Data_out <= 16'h824B	;
				14'b11000111101111: Data_out <= 16'h824E	;
				14'b11000111110000: Data_out <= 16'h8250	;
				14'b11000111110001: Data_out <= 16'h8252	;
				14'b11000111110010: Data_out <= 16'h8255	;
				14'b11000111110011: Data_out <= 16'h8257	;
				14'b11000111110100: Data_out <= 16'h825A	;
				14'b11000111110101: Data_out <= 16'h825C	;
				14'b11000111110110: Data_out <= 16'h825E	;
				14'b11000111110111: Data_out <= 16'h8261	;
				14'b11000111111000: Data_out <= 16'h8263	;
				14'b11000111111001: Data_out <= 16'h8266	;
				14'b11000111111010: Data_out <= 16'h8268	;
				14'b11000111111011: Data_out <= 16'h826B	;
				14'b11000111111100: Data_out <= 16'h826D	;
				14'b11000111111101: Data_out <= 16'h826F	;
				14'b11000111111110: Data_out <= 16'h8272	;
				14'b11000111111111: Data_out <= 16'h8274	;
				14'b11001000000000: Data_out <= 16'h8277	;
				14'b11001000000001: Data_out <= 16'h8279	;
				14'b11001000000010: Data_out <= 16'h827C	;
				14'b11001000000011: Data_out <= 16'h827E	;
				14'b11001000000100: Data_out <= 16'h8281	;
				14'b11001000000101: Data_out <= 16'h8283	;
				14'b11001000000110: Data_out <= 16'h8286	;
				14'b11001000000111: Data_out <= 16'h8288	;
				14'b11001000001000: Data_out <= 16'h828A	;
				14'b11001000001001: Data_out <= 16'h828D	;
				14'b11001000001010: Data_out <= 16'h828F	;
				14'b11001000001011: Data_out <= 16'h8292	;
				14'b11001000001100: Data_out <= 16'h8294	;
				14'b11001000001101: Data_out <= 16'h8297	;
				14'b11001000001110: Data_out <= 16'h8299	;
				14'b11001000001111: Data_out <= 16'h829C	;
				14'b11001000010000: Data_out <= 16'h829F	;
				14'b11001000010001: Data_out <= 16'h82A1	;
				14'b11001000010010: Data_out <= 16'h82A4	;
				14'b11001000010011: Data_out <= 16'h82A6	;
				14'b11001000010100: Data_out <= 16'h82A9	;
				14'b11001000010101: Data_out <= 16'h82AB	;
				14'b11001000010110: Data_out <= 16'h82AE	;
				14'b11001000010111: Data_out <= 16'h82B0	;
				14'b11001000011000: Data_out <= 16'h82B3	;
				14'b11001000011001: Data_out <= 16'h82B5	;
				14'b11001000011010: Data_out <= 16'h82B8	;
				14'b11001000011011: Data_out <= 16'h82BB	;
				14'b11001000011100: Data_out <= 16'h82BD	;
				14'b11001000011101: Data_out <= 16'h82C0	;
				14'b11001000011110: Data_out <= 16'h82C2	;
				14'b11001000011111: Data_out <= 16'h82C5	;
				14'b11001000100000: Data_out <= 16'h82C8	;
				14'b11001000100001: Data_out <= 16'h82CA	;
				14'b11001000100010: Data_out <= 16'h82CD	;
				14'b11001000100011: Data_out <= 16'h82CF	;
				14'b11001000100100: Data_out <= 16'h82D2	;
				14'b11001000100101: Data_out <= 16'h82D5	;
				14'b11001000100110: Data_out <= 16'h82D7	;
				14'b11001000100111: Data_out <= 16'h82DA	;
				14'b11001000101000: Data_out <= 16'h82DD	;
				14'b11001000101001: Data_out <= 16'h82DF	;
				14'b11001000101010: Data_out <= 16'h82E2	;
				14'b11001000101011: Data_out <= 16'h82E4	;
				14'b11001000101100: Data_out <= 16'h82E7	;
				14'b11001000101101: Data_out <= 16'h82EA	;
				14'b11001000101110: Data_out <= 16'h82EC	;
				14'b11001000101111: Data_out <= 16'h82EF	;
				14'b11001000110000: Data_out <= 16'h82F2	;
				14'b11001000110001: Data_out <= 16'h82F4	;
				14'b11001000110010: Data_out <= 16'h82F7	;
				14'b11001000110011: Data_out <= 16'h82FA	;
				14'b11001000110100: Data_out <= 16'h82FD	;
				14'b11001000110101: Data_out <= 16'h82FF	;
				14'b11001000110110: Data_out <= 16'h8302	;
				14'b11001000110111: Data_out <= 16'h8305	;
				14'b11001000111000: Data_out <= 16'h8307	;
				14'b11001000111001: Data_out <= 16'h830A	;
				14'b11001000111010: Data_out <= 16'h830D	;
				14'b11001000111011: Data_out <= 16'h8310	;
				14'b11001000111100: Data_out <= 16'h8312	;
				14'b11001000111101: Data_out <= 16'h8315	;
				14'b11001000111110: Data_out <= 16'h8318	;
				14'b11001000111111: Data_out <= 16'h831B	;
				14'b11001001000000: Data_out <= 16'h831D	;
				14'b11001001000001: Data_out <= 16'h8320	;
				14'b11001001000010: Data_out <= 16'h8323	;
				14'b11001001000011: Data_out <= 16'h8326	;
				14'b11001001000100: Data_out <= 16'h8328	;
				14'b11001001000101: Data_out <= 16'h832B	;
				14'b11001001000110: Data_out <= 16'h832E	;
				14'b11001001000111: Data_out <= 16'h8331	;
				14'b11001001001000: Data_out <= 16'h8333	;
				14'b11001001001001: Data_out <= 16'h8336	;
				14'b11001001001010: Data_out <= 16'h8339	;
				14'b11001001001011: Data_out <= 16'h833C	;
				14'b11001001001100: Data_out <= 16'h833F	;
				14'b11001001001101: Data_out <= 16'h8341	;
				14'b11001001001110: Data_out <= 16'h8344	;
				14'b11001001001111: Data_out <= 16'h8347	;
				14'b11001001010000: Data_out <= 16'h834A	;
				14'b11001001010001: Data_out <= 16'h834D	;
				14'b11001001010010: Data_out <= 16'h8350	;
				14'b11001001010011: Data_out <= 16'h8352	;
				14'b11001001010100: Data_out <= 16'h8355	;
				14'b11001001010101: Data_out <= 16'h8358	;
				14'b11001001010110: Data_out <= 16'h835B	;
				14'b11001001010111: Data_out <= 16'h835E	;
				14'b11001001011000: Data_out <= 16'h8361	;
				14'b11001001011001: Data_out <= 16'h8364	;
				14'b11001001011010: Data_out <= 16'h8366	;
				14'b11001001011011: Data_out <= 16'h8369	;
				14'b11001001011100: Data_out <= 16'h836C	;
				14'b11001001011101: Data_out <= 16'h836F	;
				14'b11001001011110: Data_out <= 16'h8372	;
				14'b11001001011111: Data_out <= 16'h8375	;
				14'b11001001100000: Data_out <= 16'h8378	;
				14'b11001001100001: Data_out <= 16'h837B	;
				14'b11001001100010: Data_out <= 16'h837E	;
				14'b11001001100011: Data_out <= 16'h8381	;
				14'b11001001100100: Data_out <= 16'h8383	;
				14'b11001001100101: Data_out <= 16'h8386	;
				14'b11001001100110: Data_out <= 16'h8389	;
				14'b11001001100111: Data_out <= 16'h838C	;
				14'b11001001101000: Data_out <= 16'h838F	;
				14'b11001001101001: Data_out <= 16'h8392	;
				14'b11001001101010: Data_out <= 16'h8395	;
				14'b11001001101011: Data_out <= 16'h8398	;
				14'b11001001101100: Data_out <= 16'h839B	;
				14'b11001001101101: Data_out <= 16'h839E	;
				14'b11001001101110: Data_out <= 16'h83A1	;
				14'b11001001101111: Data_out <= 16'h83A4	;
				14'b11001001110000: Data_out <= 16'h83A7	;
				14'b11001001110001: Data_out <= 16'h83AA	;
				14'b11001001110010: Data_out <= 16'h83AD	;
				14'b11001001110011: Data_out <= 16'h83B0	;
				14'b11001001110100: Data_out <= 16'h83B3	;
				14'b11001001110101: Data_out <= 16'h83B6	;
				14'b11001001110110: Data_out <= 16'h83B9	;
				14'b11001001110111: Data_out <= 16'h83BC	;
				14'b11001001111000: Data_out <= 16'h83BF	;
				14'b11001001111001: Data_out <= 16'h83C2	;
				14'b11001001111010: Data_out <= 16'h83C5	;
				14'b11001001111011: Data_out <= 16'h83C8	;
				14'b11001001111100: Data_out <= 16'h83CB	;
				14'b11001001111101: Data_out <= 16'h83CE	;
				14'b11001001111110: Data_out <= 16'h83D1	;
				14'b11001001111111: Data_out <= 16'h83D4	;
				14'b11001010000000: Data_out <= 16'h83D7	;
				14'b11001010000001: Data_out <= 16'h83DA	;
				14'b11001010000010: Data_out <= 16'h83DD	;
				14'b11001010000011: Data_out <= 16'h83E0	;
				14'b11001010000100: Data_out <= 16'h83E3	;
				14'b11001010000101: Data_out <= 16'h83E6	;
				14'b11001010000110: Data_out <= 16'h83E9	;
				14'b11001010000111: Data_out <= 16'h83ED	;
				14'b11001010001000: Data_out <= 16'h83F0	;
				14'b11001010001001: Data_out <= 16'h83F3	;
				14'b11001010001010: Data_out <= 16'h83F6	;
				14'b11001010001011: Data_out <= 16'h83F9	;
				14'b11001010001100: Data_out <= 16'h83FC	;
				14'b11001010001101: Data_out <= 16'h83FF	;
				14'b11001010001110: Data_out <= 16'h8402	;
				14'b11001010001111: Data_out <= 16'h8405	;
				14'b11001010010000: Data_out <= 16'h8409	;
				14'b11001010010001: Data_out <= 16'h840C	;
				14'b11001010010010: Data_out <= 16'h840F	;
				14'b11001010010011: Data_out <= 16'h8412	;
				14'b11001010010100: Data_out <= 16'h8415	;
				14'b11001010010101: Data_out <= 16'h8418	;
				14'b11001010010110: Data_out <= 16'h841B	;
				14'b11001010010111: Data_out <= 16'h841F	;
				14'b11001010011000: Data_out <= 16'h8422	;
				14'b11001010011001: Data_out <= 16'h8425	;
				14'b11001010011010: Data_out <= 16'h8428	;
				14'b11001010011011: Data_out <= 16'h842B	;
				14'b11001010011100: Data_out <= 16'h842E	;
				14'b11001010011101: Data_out <= 16'h8432	;
				14'b11001010011110: Data_out <= 16'h8435	;
				14'b11001010011111: Data_out <= 16'h8438	;
				14'b11001010100000: Data_out <= 16'h843B	;
				14'b11001010100001: Data_out <= 16'h843E	;
				14'b11001010100010: Data_out <= 16'h8442	;
				14'b11001010100011: Data_out <= 16'h8445	;
				14'b11001010100100: Data_out <= 16'h8448	;
				14'b11001010100101: Data_out <= 16'h844B	;
				14'b11001010100110: Data_out <= 16'h844E	;
				14'b11001010100111: Data_out <= 16'h8452	;
				14'b11001010101000: Data_out <= 16'h8455	;
				14'b11001010101001: Data_out <= 16'h8458	;
				14'b11001010101010: Data_out <= 16'h845B	;
				14'b11001010101011: Data_out <= 16'h845F	;
				14'b11001010101100: Data_out <= 16'h8462	;
				14'b11001010101101: Data_out <= 16'h8465	;
				14'b11001010101110: Data_out <= 16'h8468	;
				14'b11001010101111: Data_out <= 16'h846C	;
				14'b11001010110000: Data_out <= 16'h846F	;
				14'b11001010110001: Data_out <= 16'h8472	;
				14'b11001010110010: Data_out <= 16'h8476	;
				14'b11001010110011: Data_out <= 16'h8479	;
				14'b11001010110100: Data_out <= 16'h847C	;
				14'b11001010110101: Data_out <= 16'h847F	;
				14'b11001010110110: Data_out <= 16'h8483	;
				14'b11001010110111: Data_out <= 16'h8486	;
				14'b11001010111000: Data_out <= 16'h8489	;
				14'b11001010111001: Data_out <= 16'h848D	;
				14'b11001010111010: Data_out <= 16'h8490	;
				14'b11001010111011: Data_out <= 16'h8493	;
				14'b11001010111100: Data_out <= 16'h8497	;
				14'b11001010111101: Data_out <= 16'h849A	;
				14'b11001010111110: Data_out <= 16'h849D	;
				14'b11001010111111: Data_out <= 16'h84A1	;
				14'b11001011000000: Data_out <= 16'h84A4	;
				14'b11001011000001: Data_out <= 16'h84A7	;
				14'b11001011000010: Data_out <= 16'h84AB	;
				14'b11001011000011: Data_out <= 16'h84AE	;
				14'b11001011000100: Data_out <= 16'h84B1	;
				14'b11001011000101: Data_out <= 16'h84B5	;
				14'b11001011000110: Data_out <= 16'h84B8	;
				14'b11001011000111: Data_out <= 16'h84BC	;
				14'b11001011001000: Data_out <= 16'h84BF	;
				14'b11001011001001: Data_out <= 16'h84C2	;
				14'b11001011001010: Data_out <= 16'h84C6	;
				14'b11001011001011: Data_out <= 16'h84C9	;
				14'b11001011001100: Data_out <= 16'h84CD	;
				14'b11001011001101: Data_out <= 16'h84D0	;
				14'b11001011001110: Data_out <= 16'h84D3	;
				14'b11001011001111: Data_out <= 16'h84D7	;
				14'b11001011010000: Data_out <= 16'h84DA	;
				14'b11001011010001: Data_out <= 16'h84DE	;
				14'b11001011010010: Data_out <= 16'h84E1	;
				14'b11001011010011: Data_out <= 16'h84E5	;
				14'b11001011010100: Data_out <= 16'h84E8	;
				14'b11001011010101: Data_out <= 16'h84EB	;
				14'b11001011010110: Data_out <= 16'h84EF	;
				14'b11001011010111: Data_out <= 16'h84F2	;
				14'b11001011011000: Data_out <= 16'h84F6	;
				14'b11001011011001: Data_out <= 16'h84F9	;
				14'b11001011011010: Data_out <= 16'h84FD	;
				14'b11001011011011: Data_out <= 16'h8500	;
				14'b11001011011100: Data_out <= 16'h8504	;
				14'b11001011011101: Data_out <= 16'h8507	;
				14'b11001011011110: Data_out <= 16'h850B	;
				14'b11001011011111: Data_out <= 16'h850E	;
				14'b11001011100000: Data_out <= 16'h8512	;
				14'b11001011100001: Data_out <= 16'h8515	;
				14'b11001011100010: Data_out <= 16'h8519	;
				14'b11001011100011: Data_out <= 16'h851C	;
				14'b11001011100100: Data_out <= 16'h8520	;
				14'b11001011100101: Data_out <= 16'h8523	;
				14'b11001011100110: Data_out <= 16'h8527	;
				14'b11001011100111: Data_out <= 16'h852A	;
				14'b11001011101000: Data_out <= 16'h852E	;
				14'b11001011101001: Data_out <= 16'h8531	;
				14'b11001011101010: Data_out <= 16'h8535	;
				14'b11001011101011: Data_out <= 16'h8538	;
				14'b11001011101100: Data_out <= 16'h853C	;
				14'b11001011101101: Data_out <= 16'h8540	;
				14'b11001011101110: Data_out <= 16'h8543	;
				14'b11001011101111: Data_out <= 16'h8547	;
				14'b11001011110000: Data_out <= 16'h854A	;
				14'b11001011110001: Data_out <= 16'h854E	;
				14'b11001011110010: Data_out <= 16'h8551	;
				14'b11001011110011: Data_out <= 16'h8555	;
				14'b11001011110100: Data_out <= 16'h8559	;
				14'b11001011110101: Data_out <= 16'h855C	;
				14'b11001011110110: Data_out <= 16'h8560	;
				14'b11001011110111: Data_out <= 16'h8563	;
				14'b11001011111000: Data_out <= 16'h8567	;
				14'b11001011111001: Data_out <= 16'h856B	;
				14'b11001011111010: Data_out <= 16'h856E	;
				14'b11001011111011: Data_out <= 16'h8572	;
				14'b11001011111100: Data_out <= 16'h8575	;
				14'b11001011111101: Data_out <= 16'h8579	;
				14'b11001011111110: Data_out <= 16'h857D	;
				14'b11001011111111: Data_out <= 16'h8580	;
				14'b11001100000000: Data_out <= 16'h8584	;
				14'b11001100000001: Data_out <= 16'h8588	;
				14'b11001100000010: Data_out <= 16'h858B	;
				14'b11001100000011: Data_out <= 16'h858F	;
				14'b11001100000100: Data_out <= 16'h8593	;
				14'b11001100000101: Data_out <= 16'h8596	;
				14'b11001100000110: Data_out <= 16'h859A	;
				14'b11001100000111: Data_out <= 16'h859E	;
				14'b11001100001000: Data_out <= 16'h85A1	;
				14'b11001100001001: Data_out <= 16'h85A5	;
				14'b11001100001010: Data_out <= 16'h85A9	;
				14'b11001100001011: Data_out <= 16'h85AC	;
				14'b11001100001100: Data_out <= 16'h85B0	;
				14'b11001100001101: Data_out <= 16'h85B4	;
				14'b11001100001110: Data_out <= 16'h85B8	;
				14'b11001100001111: Data_out <= 16'h85BB	;
				14'b11001100010000: Data_out <= 16'h85BF	;
				14'b11001100010001: Data_out <= 16'h85C3	;
				14'b11001100010010: Data_out <= 16'h85C6	;
				14'b11001100010011: Data_out <= 16'h85CA	;
				14'b11001100010100: Data_out <= 16'h85CE	;
				14'b11001100010101: Data_out <= 16'h85D2	;
				14'b11001100010110: Data_out <= 16'h85D5	;
				14'b11001100010111: Data_out <= 16'h85D9	;
				14'b11001100011000: Data_out <= 16'h85DD	;
				14'b11001100011001: Data_out <= 16'h85E1	;
				14'b11001100011010: Data_out <= 16'h85E4	;
				14'b11001100011011: Data_out <= 16'h85E8	;
				14'b11001100011100: Data_out <= 16'h85EC	;
				14'b11001100011101: Data_out <= 16'h85F0	;
				14'b11001100011110: Data_out <= 16'h85F4	;
				14'b11001100011111: Data_out <= 16'h85F7	;
				14'b11001100100000: Data_out <= 16'h85FB	;
				14'b11001100100001: Data_out <= 16'h85FF	;
				14'b11001100100010: Data_out <= 16'h8603	;
				14'b11001100100011: Data_out <= 16'h8607	;
				14'b11001100100100: Data_out <= 16'h860A	;
				14'b11001100100101: Data_out <= 16'h860E	;
				14'b11001100100110: Data_out <= 16'h8612	;
				14'b11001100100111: Data_out <= 16'h8616	;
				14'b11001100101000: Data_out <= 16'h861A	;
				14'b11001100101001: Data_out <= 16'h861D	;
				14'b11001100101010: Data_out <= 16'h8621	;
				14'b11001100101011: Data_out <= 16'h8625	;
				14'b11001100101100: Data_out <= 16'h8629	;
				14'b11001100101101: Data_out <= 16'h862D	;
				14'b11001100101110: Data_out <= 16'h8631	;
				14'b11001100101111: Data_out <= 16'h8635	;
				14'b11001100110000: Data_out <= 16'h8638	;
				14'b11001100110001: Data_out <= 16'h863C	;
				14'b11001100110010: Data_out <= 16'h8640	;
				14'b11001100110011: Data_out <= 16'h8644	;
				14'b11001100110100: Data_out <= 16'h8648	;
				14'b11001100110101: Data_out <= 16'h864C	;
				14'b11001100110110: Data_out <= 16'h8650	;
				14'b11001100110111: Data_out <= 16'h8654	;
				14'b11001100111000: Data_out <= 16'h8658	;
				14'b11001100111001: Data_out <= 16'h865B	;
				14'b11001100111010: Data_out <= 16'h865F	;
				14'b11001100111011: Data_out <= 16'h8663	;
				14'b11001100111100: Data_out <= 16'h8667	;
				14'b11001100111101: Data_out <= 16'h866B	;
				14'b11001100111110: Data_out <= 16'h866F	;
				14'b11001100111111: Data_out <= 16'h8673	;
				14'b11001101000000: Data_out <= 16'h8677	;
				14'b11001101000001: Data_out <= 16'h867B	;
				14'b11001101000010: Data_out <= 16'h867F	;
				14'b11001101000011: Data_out <= 16'h8683	;
				14'b11001101000100: Data_out <= 16'h8687	;
				14'b11001101000101: Data_out <= 16'h868B	;
				14'b11001101000110: Data_out <= 16'h868F	;
				14'b11001101000111: Data_out <= 16'h8693	;
				14'b11001101001000: Data_out <= 16'h8697	;
				14'b11001101001001: Data_out <= 16'h869B	;
				14'b11001101001010: Data_out <= 16'h869F	;
				14'b11001101001011: Data_out <= 16'h86A3	;
				14'b11001101001100: Data_out <= 16'h86A7	;
				14'b11001101001101: Data_out <= 16'h86AB	;
				14'b11001101001110: Data_out <= 16'h86AF	;
				14'b11001101001111: Data_out <= 16'h86B3	;
				14'b11001101010000: Data_out <= 16'h86B7	;
				14'b11001101010001: Data_out <= 16'h86BB	;
				14'b11001101010010: Data_out <= 16'h86BF	;
				14'b11001101010011: Data_out <= 16'h86C3	;
				14'b11001101010100: Data_out <= 16'h86C7	;
				14'b11001101010101: Data_out <= 16'h86CB	;
				14'b11001101010110: Data_out <= 16'h86CF	;
				14'b11001101010111: Data_out <= 16'h86D3	;
				14'b11001101011000: Data_out <= 16'h86D7	;
				14'b11001101011001: Data_out <= 16'h86DB	;
				14'b11001101011010: Data_out <= 16'h86DF	;
				14'b11001101011011: Data_out <= 16'h86E3	;
				14'b11001101011100: Data_out <= 16'h86E7	;
				14'b11001101011101: Data_out <= 16'h86EB	;
				14'b11001101011110: Data_out <= 16'h86EF	;
				14'b11001101011111: Data_out <= 16'h86F3	;
				14'b11001101100000: Data_out <= 16'h86F7	;
				14'b11001101100001: Data_out <= 16'h86FB	;
				14'b11001101100010: Data_out <= 16'h8700	;
				14'b11001101100011: Data_out <= 16'h8704	;
				14'b11001101100100: Data_out <= 16'h8708	;
				14'b11001101100101: Data_out <= 16'h870C	;
				14'b11001101100110: Data_out <= 16'h8710	;
				14'b11001101100111: Data_out <= 16'h8714	;
				14'b11001101101000: Data_out <= 16'h8718	;
				14'b11001101101001: Data_out <= 16'h871C	;
				14'b11001101101010: Data_out <= 16'h8720	;
				14'b11001101101011: Data_out <= 16'h8725	;
				14'b11001101101100: Data_out <= 16'h8729	;
				14'b11001101101101: Data_out <= 16'h872D	;
				14'b11001101101110: Data_out <= 16'h8731	;
				14'b11001101101111: Data_out <= 16'h8735	;
				14'b11001101110000: Data_out <= 16'h8739	;
				14'b11001101110001: Data_out <= 16'h873E	;
				14'b11001101110010: Data_out <= 16'h8742	;
				14'b11001101110011: Data_out <= 16'h8746	;
				14'b11001101110100: Data_out <= 16'h874A	;
				14'b11001101110101: Data_out <= 16'h874E	;
				14'b11001101110110: Data_out <= 16'h8752	;
				14'b11001101110111: Data_out <= 16'h8757	;
				14'b11001101111000: Data_out <= 16'h875B	;
				14'b11001101111001: Data_out <= 16'h875F	;
				14'b11001101111010: Data_out <= 16'h8763	;
				14'b11001101111011: Data_out <= 16'h8767	;
				14'b11001101111100: Data_out <= 16'h876C	;
				14'b11001101111101: Data_out <= 16'h8770	;
				14'b11001101111110: Data_out <= 16'h8774	;
				14'b11001101111111: Data_out <= 16'h8778	;
				14'b11001110000000: Data_out <= 16'h877D	;
				14'b11001110000001: Data_out <= 16'h8781	;
				14'b11001110000010: Data_out <= 16'h8785	;
				14'b11001110000011: Data_out <= 16'h8789	;
				14'b11001110000100: Data_out <= 16'h878D	;
				14'b11001110000101: Data_out <= 16'h8792	;
				14'b11001110000110: Data_out <= 16'h8796	;
				14'b11001110000111: Data_out <= 16'h879A	;
				14'b11001110001000: Data_out <= 16'h879F	;
				14'b11001110001001: Data_out <= 16'h87A3	;
				14'b11001110001010: Data_out <= 16'h87A7	;
				14'b11001110001011: Data_out <= 16'h87AB	;
				14'b11001110001100: Data_out <= 16'h87B0	;
				14'b11001110001101: Data_out <= 16'h87B4	;
				14'b11001110001110: Data_out <= 16'h87B8	;
				14'b11001110001111: Data_out <= 16'h87BD	;
				14'b11001110010000: Data_out <= 16'h87C1	;
				14'b11001110010001: Data_out <= 16'h87C5	;
				14'b11001110010010: Data_out <= 16'h87C9	;
				14'b11001110010011: Data_out <= 16'h87CE	;
				14'b11001110010100: Data_out <= 16'h87D2	;
				14'b11001110010101: Data_out <= 16'h87D6	;
				14'b11001110010110: Data_out <= 16'h87DB	;
				14'b11001110010111: Data_out <= 16'h87DF	;
				14'b11001110011000: Data_out <= 16'h87E3	;
				14'b11001110011001: Data_out <= 16'h87E8	;
				14'b11001110011010: Data_out <= 16'h87EC	;
				14'b11001110011011: Data_out <= 16'h87F0	;
				14'b11001110011100: Data_out <= 16'h87F5	;
				14'b11001110011101: Data_out <= 16'h87F9	;
				14'b11001110011110: Data_out <= 16'h87FE	;
				14'b11001110011111: Data_out <= 16'h8802	;
				14'b11001110100000: Data_out <= 16'h8806	;
				14'b11001110100001: Data_out <= 16'h880B	;
				14'b11001110100010: Data_out <= 16'h880F	;
				14'b11001110100011: Data_out <= 16'h8813	;
				14'b11001110100100: Data_out <= 16'h8818	;
				14'b11001110100101: Data_out <= 16'h881C	;
				14'b11001110100110: Data_out <= 16'h8821	;
				14'b11001110100111: Data_out <= 16'h8825	;
				14'b11001110101000: Data_out <= 16'h8829	;
				14'b11001110101001: Data_out <= 16'h882E	;
				14'b11001110101010: Data_out <= 16'h8832	;
				14'b11001110101011: Data_out <= 16'h8837	;
				14'b11001110101100: Data_out <= 16'h883B	;
				14'b11001110101101: Data_out <= 16'h8840	;
				14'b11001110101110: Data_out <= 16'h8844	;
				14'b11001110101111: Data_out <= 16'h8848	;
				14'b11001110110000: Data_out <= 16'h884D	;
				14'b11001110110001: Data_out <= 16'h8851	;
				14'b11001110110010: Data_out <= 16'h8856	;
				14'b11001110110011: Data_out <= 16'h885A	;
				14'b11001110110100: Data_out <= 16'h885F	;
				14'b11001110110101: Data_out <= 16'h8863	;
				14'b11001110110110: Data_out <= 16'h8868	;
				14'b11001110110111: Data_out <= 16'h886C	;
				14'b11001110111000: Data_out <= 16'h8871	;
				14'b11001110111001: Data_out <= 16'h8875	;
				14'b11001110111010: Data_out <= 16'h887A	;
				14'b11001110111011: Data_out <= 16'h887E	;
				14'b11001110111100: Data_out <= 16'h8883	;
				14'b11001110111101: Data_out <= 16'h8887	;
				14'b11001110111110: Data_out <= 16'h888C	;
				14'b11001110111111: Data_out <= 16'h8890	;
				14'b11001111000000: Data_out <= 16'h8895	;
				14'b11001111000001: Data_out <= 16'h8899	;
				14'b11001111000010: Data_out <= 16'h889E	;
				14'b11001111000011: Data_out <= 16'h88A2	;
				14'b11001111000100: Data_out <= 16'h88A7	;
				14'b11001111000101: Data_out <= 16'h88AB	;
				14'b11001111000110: Data_out <= 16'h88B0	;
				14'b11001111000111: Data_out <= 16'h88B4	;
				14'b11001111001000: Data_out <= 16'h88B9	;
				14'b11001111001001: Data_out <= 16'h88BE	;
				14'b11001111001010: Data_out <= 16'h88C2	;
				14'b11001111001011: Data_out <= 16'h88C7	;
				14'b11001111001100: Data_out <= 16'h88CB	;
				14'b11001111001101: Data_out <= 16'h88D0	;
				14'b11001111001110: Data_out <= 16'h88D4	;
				14'b11001111001111: Data_out <= 16'h88D9	;
				14'b11001111010000: Data_out <= 16'h88DE	;
				14'b11001111010001: Data_out <= 16'h88E2	;
				14'b11001111010010: Data_out <= 16'h88E7	;
				14'b11001111010011: Data_out <= 16'h88EB	;
				14'b11001111010100: Data_out <= 16'h88F0	;
				14'b11001111010101: Data_out <= 16'h88F5	;
				14'b11001111010110: Data_out <= 16'h88F9	;
				14'b11001111010111: Data_out <= 16'h88FE	;
				14'b11001111011000: Data_out <= 16'h8903	;
				14'b11001111011001: Data_out <= 16'h8907	;
				14'b11001111011010: Data_out <= 16'h890C	;
				14'b11001111011011: Data_out <= 16'h8910	;
				14'b11001111011100: Data_out <= 16'h8915	;
				14'b11001111011101: Data_out <= 16'h891A	;
				14'b11001111011110: Data_out <= 16'h891E	;
				14'b11001111011111: Data_out <= 16'h8923	;
				14'b11001111100000: Data_out <= 16'h8928	;
				14'b11001111100001: Data_out <= 16'h892C	;
				14'b11001111100010: Data_out <= 16'h8931	;
				14'b11001111100011: Data_out <= 16'h8936	;
				14'b11001111100100: Data_out <= 16'h893A	;
				14'b11001111100101: Data_out <= 16'h893F	;
				14'b11001111100110: Data_out <= 16'h8944	;
				14'b11001111100111: Data_out <= 16'h8949	;
				14'b11001111101000: Data_out <= 16'h894D	;
				14'b11001111101001: Data_out <= 16'h8952	;
				14'b11001111101010: Data_out <= 16'h8957	;
				14'b11001111101011: Data_out <= 16'h895B	;
				14'b11001111101100: Data_out <= 16'h8960	;
				14'b11001111101101: Data_out <= 16'h8965	;
				14'b11001111101110: Data_out <= 16'h896A	;
				14'b11001111101111: Data_out <= 16'h896E	;
				14'b11001111110000: Data_out <= 16'h8973	;
				14'b11001111110001: Data_out <= 16'h8978	;
				14'b11001111110010: Data_out <= 16'h897C	;
				14'b11001111110011: Data_out <= 16'h8981	;
				14'b11001111110100: Data_out <= 16'h8986	;
				14'b11001111110101: Data_out <= 16'h898B	;
				14'b11001111110110: Data_out <= 16'h898F	;
				14'b11001111110111: Data_out <= 16'h8994	;
				14'b11001111111000: Data_out <= 16'h8999	;
				14'b11001111111001: Data_out <= 16'h899E	;
				14'b11001111111010: Data_out <= 16'h89A3	;
				14'b11001111111011: Data_out <= 16'h89A7	;
				14'b11001111111100: Data_out <= 16'h89AC	;
				14'b11001111111101: Data_out <= 16'h89B1	;
				14'b11001111111110: Data_out <= 16'h89B6	;
				14'b11001111111111: Data_out <= 16'h89BB	;
				14'b11010000000000: Data_out <= 16'h89BF	;
				14'b11010000000001: Data_out <= 16'h89C4	;
				14'b11010000000010: Data_out <= 16'h89C9	;
				14'b11010000000011: Data_out <= 16'h89CE	;
				14'b11010000000100: Data_out <= 16'h89D3	;
				14'b11010000000101: Data_out <= 16'h89D7	;
				14'b11010000000110: Data_out <= 16'h89DC	;
				14'b11010000000111: Data_out <= 16'h89E1	;
				14'b11010000001000: Data_out <= 16'h89E6	;
				14'b11010000001001: Data_out <= 16'h89EB	;
				14'b11010000001010: Data_out <= 16'h89F0	;
				14'b11010000001011: Data_out <= 16'h89F5	;
				14'b11010000001100: Data_out <= 16'h89F9	;
				14'b11010000001101: Data_out <= 16'h89FE	;
				14'b11010000001110: Data_out <= 16'h8A03	;
				14'b11010000001111: Data_out <= 16'h8A08	;
				14'b11010000010000: Data_out <= 16'h8A0D	;
				14'b11010000010001: Data_out <= 16'h8A12	;
				14'b11010000010010: Data_out <= 16'h8A17	;
				14'b11010000010011: Data_out <= 16'h8A1C	;
				14'b11010000010100: Data_out <= 16'h8A20	;
				14'b11010000010101: Data_out <= 16'h8A25	;
				14'b11010000010110: Data_out <= 16'h8A2A	;
				14'b11010000010111: Data_out <= 16'h8A2F	;
				14'b11010000011000: Data_out <= 16'h8A34	;
				14'b11010000011001: Data_out <= 16'h8A39	;
				14'b11010000011010: Data_out <= 16'h8A3E	;
				14'b11010000011011: Data_out <= 16'h8A43	;
				14'b11010000011100: Data_out <= 16'h8A48	;
				14'b11010000011101: Data_out <= 16'h8A4D	;
				14'b11010000011110: Data_out <= 16'h8A52	;
				14'b11010000011111: Data_out <= 16'h8A57	;
				14'b11010000100000: Data_out <= 16'h8A5B	;
				14'b11010000100001: Data_out <= 16'h8A60	;
				14'b11010000100010: Data_out <= 16'h8A65	;
				14'b11010000100011: Data_out <= 16'h8A6A	;
				14'b11010000100100: Data_out <= 16'h8A6F	;
				14'b11010000100101: Data_out <= 16'h8A74	;
				14'b11010000100110: Data_out <= 16'h8A79	;
				14'b11010000100111: Data_out <= 16'h8A7E	;
				14'b11010000101000: Data_out <= 16'h8A83	;
				14'b11010000101001: Data_out <= 16'h8A88	;
				14'b11010000101010: Data_out <= 16'h8A8D	;
				14'b11010000101011: Data_out <= 16'h8A92	;
				14'b11010000101100: Data_out <= 16'h8A97	;
				14'b11010000101101: Data_out <= 16'h8A9C	;
				14'b11010000101110: Data_out <= 16'h8AA1	;
				14'b11010000101111: Data_out <= 16'h8AA6	;
				14'b11010000110000: Data_out <= 16'h8AAB	;
				14'b11010000110001: Data_out <= 16'h8AB0	;
				14'b11010000110010: Data_out <= 16'h8AB5	;
				14'b11010000110011: Data_out <= 16'h8ABA	;
				14'b11010000110100: Data_out <= 16'h8ABF	;
				14'b11010000110101: Data_out <= 16'h8AC4	;
				14'b11010000110110: Data_out <= 16'h8AC9	;
				14'b11010000110111: Data_out <= 16'h8ACF	;
				14'b11010000111000: Data_out <= 16'h8AD4	;
				14'b11010000111001: Data_out <= 16'h8AD9	;
				14'b11010000111010: Data_out <= 16'h8ADE	;
				14'b11010000111011: Data_out <= 16'h8AE3	;
				14'b11010000111100: Data_out <= 16'h8AE8	;
				14'b11010000111101: Data_out <= 16'h8AED	;
				14'b11010000111110: Data_out <= 16'h8AF2	;
				14'b11010000111111: Data_out <= 16'h8AF7	;
				14'b11010001000000: Data_out <= 16'h8AFC	;
				14'b11010001000001: Data_out <= 16'h8B01	;
				14'b11010001000010: Data_out <= 16'h8B06	;
				14'b11010001000011: Data_out <= 16'h8B0B	;
				14'b11010001000100: Data_out <= 16'h8B11	;
				14'b11010001000101: Data_out <= 16'h8B16	;
				14'b11010001000110: Data_out <= 16'h8B1B	;
				14'b11010001000111: Data_out <= 16'h8B20	;
				14'b11010001001000: Data_out <= 16'h8B25	;
				14'b11010001001001: Data_out <= 16'h8B2A	;
				14'b11010001001010: Data_out <= 16'h8B2F	;
				14'b11010001001011: Data_out <= 16'h8B34	;
				14'b11010001001100: Data_out <= 16'h8B3A	;
				14'b11010001001101: Data_out <= 16'h8B3F	;
				14'b11010001001110: Data_out <= 16'h8B44	;
				14'b11010001001111: Data_out <= 16'h8B49	;
				14'b11010001010000: Data_out <= 16'h8B4E	;
				14'b11010001010001: Data_out <= 16'h8B53	;
				14'b11010001010010: Data_out <= 16'h8B59	;
				14'b11010001010011: Data_out <= 16'h8B5E	;
				14'b11010001010100: Data_out <= 16'h8B63	;
				14'b11010001010101: Data_out <= 16'h8B68	;
				14'b11010001010110: Data_out <= 16'h8B6D	;
				14'b11010001010111: Data_out <= 16'h8B72	;
				14'b11010001011000: Data_out <= 16'h8B78	;
				14'b11010001011001: Data_out <= 16'h8B7D	;
				14'b11010001011010: Data_out <= 16'h8B82	;
				14'b11010001011011: Data_out <= 16'h8B87	;
				14'b11010001011100: Data_out <= 16'h8B8C	;
				14'b11010001011101: Data_out <= 16'h8B92	;
				14'b11010001011110: Data_out <= 16'h8B97	;
				14'b11010001011111: Data_out <= 16'h8B9C	;
				14'b11010001100000: Data_out <= 16'h8BA1	;
				14'b11010001100001: Data_out <= 16'h8BA7	;
				14'b11010001100010: Data_out <= 16'h8BAC	;
				14'b11010001100011: Data_out <= 16'h8BB1	;
				14'b11010001100100: Data_out <= 16'h8BB6	;
				14'b11010001100101: Data_out <= 16'h8BBC	;
				14'b11010001100110: Data_out <= 16'h8BC1	;
				14'b11010001100111: Data_out <= 16'h8BC6	;
				14'b11010001101000: Data_out <= 16'h8BCB	;
				14'b11010001101001: Data_out <= 16'h8BD1	;
				14'b11010001101010: Data_out <= 16'h8BD6	;
				14'b11010001101011: Data_out <= 16'h8BDB	;
				14'b11010001101100: Data_out <= 16'h8BE1	;
				14'b11010001101101: Data_out <= 16'h8BE6	;
				14'b11010001101110: Data_out <= 16'h8BEB	;
				14'b11010001101111: Data_out <= 16'h8BF0	;
				14'b11010001110000: Data_out <= 16'h8BF6	;
				14'b11010001110001: Data_out <= 16'h8BFB	;
				14'b11010001110010: Data_out <= 16'h8C00	;
				14'b11010001110011: Data_out <= 16'h8C06	;
				14'b11010001110100: Data_out <= 16'h8C0B	;
				14'b11010001110101: Data_out <= 16'h8C10	;
				14'b11010001110110: Data_out <= 16'h8C16	;
				14'b11010001110111: Data_out <= 16'h8C1B	;
				14'b11010001111000: Data_out <= 16'h8C20	;
				14'b11010001111001: Data_out <= 16'h8C26	;
				14'b11010001111010: Data_out <= 16'h8C2B	;
				14'b11010001111011: Data_out <= 16'h8C30	;
				14'b11010001111100: Data_out <= 16'h8C36	;
				14'b11010001111101: Data_out <= 16'h8C3B	;
				14'b11010001111110: Data_out <= 16'h8C40	;
				14'b11010001111111: Data_out <= 16'h8C46	;
				14'b11010010000000: Data_out <= 16'h8C4B	;
				14'b11010010000001: Data_out <= 16'h8C50	;
				14'b11010010000010: Data_out <= 16'h8C56	;
				14'b11010010000011: Data_out <= 16'h8C5B	;
				14'b11010010000100: Data_out <= 16'h8C61	;
				14'b11010010000101: Data_out <= 16'h8C66	;
				14'b11010010000110: Data_out <= 16'h8C6B	;
				14'b11010010000111: Data_out <= 16'h8C71	;
				14'b11010010001000: Data_out <= 16'h8C76	;
				14'b11010010001001: Data_out <= 16'h8C7C	;
				14'b11010010001010: Data_out <= 16'h8C81	;
				14'b11010010001011: Data_out <= 16'h8C86	;
				14'b11010010001100: Data_out <= 16'h8C8C	;
				14'b11010010001101: Data_out <= 16'h8C91	;
				14'b11010010001110: Data_out <= 16'h8C97	;
				14'b11010010001111: Data_out <= 16'h8C9C	;
				14'b11010010010000: Data_out <= 16'h8CA2	;
				14'b11010010010001: Data_out <= 16'h8CA7	;
				14'b11010010010010: Data_out <= 16'h8CAC	;
				14'b11010010010011: Data_out <= 16'h8CB2	;
				14'b11010010010100: Data_out <= 16'h8CB7	;
				14'b11010010010101: Data_out <= 16'h8CBD	;
				14'b11010010010110: Data_out <= 16'h8CC2	;
				14'b11010010010111: Data_out <= 16'h8CC8	;
				14'b11010010011000: Data_out <= 16'h8CCD	;
				14'b11010010011001: Data_out <= 16'h8CD3	;
				14'b11010010011010: Data_out <= 16'h8CD8	;
				14'b11010010011011: Data_out <= 16'h8CDE	;
				14'b11010010011100: Data_out <= 16'h8CE3	;
				14'b11010010011101: Data_out <= 16'h8CE9	;
				14'b11010010011110: Data_out <= 16'h8CEE	;
				14'b11010010011111: Data_out <= 16'h8CF4	;
				14'b11010010100000: Data_out <= 16'h8CF9	;
				14'b11010010100001: Data_out <= 16'h8CFF	;
				14'b11010010100010: Data_out <= 16'h8D04	;
				14'b11010010100011: Data_out <= 16'h8D0A	;
				14'b11010010100100: Data_out <= 16'h8D0F	;
				14'b11010010100101: Data_out <= 16'h8D15	;
				14'b11010010100110: Data_out <= 16'h8D1A	;
				14'b11010010100111: Data_out <= 16'h8D20	;
				14'b11010010101000: Data_out <= 16'h8D25	;
				14'b11010010101001: Data_out <= 16'h8D2B	;
				14'b11010010101010: Data_out <= 16'h8D31	;
				14'b11010010101011: Data_out <= 16'h8D36	;
				14'b11010010101100: Data_out <= 16'h8D3C	;
				14'b11010010101101: Data_out <= 16'h8D41	;
				14'b11010010101110: Data_out <= 16'h8D47	;
				14'b11010010101111: Data_out <= 16'h8D4C	;
				14'b11010010110000: Data_out <= 16'h8D52	;
				14'b11010010110001: Data_out <= 16'h8D58	;
				14'b11010010110010: Data_out <= 16'h8D5D	;
				14'b11010010110011: Data_out <= 16'h8D63	;
				14'b11010010110100: Data_out <= 16'h8D68	;
				14'b11010010110101: Data_out <= 16'h8D6E	;
				14'b11010010110110: Data_out <= 16'h8D74	;
				14'b11010010110111: Data_out <= 16'h8D79	;
				14'b11010010111000: Data_out <= 16'h8D7F	;
				14'b11010010111001: Data_out <= 16'h8D84	;
				14'b11010010111010: Data_out <= 16'h8D8A	;
				14'b11010010111011: Data_out <= 16'h8D90	;
				14'b11010010111100: Data_out <= 16'h8D95	;
				14'b11010010111101: Data_out <= 16'h8D9B	;
				14'b11010010111110: Data_out <= 16'h8DA1	;
				14'b11010010111111: Data_out <= 16'h8DA6	;
				14'b11010011000000: Data_out <= 16'h8DAC	;
				14'b11010011000001: Data_out <= 16'h8DB1	;
				14'b11010011000010: Data_out <= 16'h8DB7	;
				14'b11010011000011: Data_out <= 16'h8DBD	;
				14'b11010011000100: Data_out <= 16'h8DC2	;
				14'b11010011000101: Data_out <= 16'h8DC8	;
				14'b11010011000110: Data_out <= 16'h8DCE	;
				14'b11010011000111: Data_out <= 16'h8DD3	;
				14'b11010011001000: Data_out <= 16'h8DD9	;
				14'b11010011001001: Data_out <= 16'h8DDF	;
				14'b11010011001010: Data_out <= 16'h8DE5	;
				14'b11010011001011: Data_out <= 16'h8DEA	;
				14'b11010011001100: Data_out <= 16'h8DF0	;
				14'b11010011001101: Data_out <= 16'h8DF6	;
				14'b11010011001110: Data_out <= 16'h8DFB	;
				14'b11010011001111: Data_out <= 16'h8E01	;
				14'b11010011010000: Data_out <= 16'h8E07	;
				14'b11010011010001: Data_out <= 16'h8E0C	;
				14'b11010011010010: Data_out <= 16'h8E12	;
				14'b11010011010011: Data_out <= 16'h8E18	;
				14'b11010011010100: Data_out <= 16'h8E1E	;
				14'b11010011010101: Data_out <= 16'h8E23	;
				14'b11010011010110: Data_out <= 16'h8E29	;
				14'b11010011010111: Data_out <= 16'h8E2F	;
				14'b11010011011000: Data_out <= 16'h8E35	;
				14'b11010011011001: Data_out <= 16'h8E3A	;
				14'b11010011011010: Data_out <= 16'h8E40	;
				14'b11010011011011: Data_out <= 16'h8E46	;
				14'b11010011011100: Data_out <= 16'h8E4C	;
				14'b11010011011101: Data_out <= 16'h8E51	;
				14'b11010011011110: Data_out <= 16'h8E57	;
				14'b11010011011111: Data_out <= 16'h8E5D	;
				14'b11010011100000: Data_out <= 16'h8E63	;
				14'b11010011100001: Data_out <= 16'h8E69	;
				14'b11010011100010: Data_out <= 16'h8E6E	;
				14'b11010011100011: Data_out <= 16'h8E74	;
				14'b11010011100100: Data_out <= 16'h8E7A	;
				14'b11010011100101: Data_out <= 16'h8E80	;
				14'b11010011100110: Data_out <= 16'h8E86	;
				14'b11010011100111: Data_out <= 16'h8E8B	;
				14'b11010011101000: Data_out <= 16'h8E91	;
				14'b11010011101001: Data_out <= 16'h8E97	;
				14'b11010011101010: Data_out <= 16'h8E9D	;
				14'b11010011101011: Data_out <= 16'h8EA3	;
				14'b11010011101100: Data_out <= 16'h8EA9	;
				14'b11010011101101: Data_out <= 16'h8EAE	;
				14'b11010011101110: Data_out <= 16'h8EB4	;
				14'b11010011101111: Data_out <= 16'h8EBA	;
				14'b11010011110000: Data_out <= 16'h8EC0	;
				14'b11010011110001: Data_out <= 16'h8EC6	;
				14'b11010011110010: Data_out <= 16'h8ECC	;
				14'b11010011110011: Data_out <= 16'h8ED2	;
				14'b11010011110100: Data_out <= 16'h8ED7	;
				14'b11010011110101: Data_out <= 16'h8EDD	;
				14'b11010011110110: Data_out <= 16'h8EE3	;
				14'b11010011110111: Data_out <= 16'h8EE9	;
				14'b11010011111000: Data_out <= 16'h8EEF	;
				14'b11010011111001: Data_out <= 16'h8EF5	;
				14'b11010011111010: Data_out <= 16'h8EFB	;
				14'b11010011111011: Data_out <= 16'h8F01	;
				14'b11010011111100: Data_out <= 16'h8F07	;
				14'b11010011111101: Data_out <= 16'h8F0C	;
				14'b11010011111110: Data_out <= 16'h8F12	;
				14'b11010011111111: Data_out <= 16'h8F18	;
				14'b11010100000000: Data_out <= 16'h8F1E	;
				14'b11010100000001: Data_out <= 16'h8F24	;
				14'b11010100000010: Data_out <= 16'h8F2A	;
				14'b11010100000011: Data_out <= 16'h8F30	;
				14'b11010100000100: Data_out <= 16'h8F36	;
				14'b11010100000101: Data_out <= 16'h8F3C	;
				14'b11010100000110: Data_out <= 16'h8F42	;
				14'b11010100000111: Data_out <= 16'h8F48	;
				14'b11010100001000: Data_out <= 16'h8F4E	;
				14'b11010100001001: Data_out <= 16'h8F54	;
				14'b11010100001010: Data_out <= 16'h8F5A	;
				14'b11010100001011: Data_out <= 16'h8F60	;
				14'b11010100001100: Data_out <= 16'h8F66	;
				14'b11010100001101: Data_out <= 16'h8F6C	;
				14'b11010100001110: Data_out <= 16'h8F72	;
				14'b11010100001111: Data_out <= 16'h8F78	;
				14'b11010100010000: Data_out <= 16'h8F7E	;
				14'b11010100010001: Data_out <= 16'h8F83	;
				14'b11010100010010: Data_out <= 16'h8F89	;
				14'b11010100010011: Data_out <= 16'h8F8F	;
				14'b11010100010100: Data_out <= 16'h8F96	;
				14'b11010100010101: Data_out <= 16'h8F9C	;
				14'b11010100010110: Data_out <= 16'h8FA2	;
				14'b11010100010111: Data_out <= 16'h8FA8	;
				14'b11010100011000: Data_out <= 16'h8FAE	;
				14'b11010100011001: Data_out <= 16'h8FB4	;
				14'b11010100011010: Data_out <= 16'h8FBA	;
				14'b11010100011011: Data_out <= 16'h8FC0	;
				14'b11010100011100: Data_out <= 16'h8FC6	;
				14'b11010100011101: Data_out <= 16'h8FCC	;
				14'b11010100011110: Data_out <= 16'h8FD2	;
				14'b11010100011111: Data_out <= 16'h8FD8	;
				14'b11010100100000: Data_out <= 16'h8FDE	;
				14'b11010100100001: Data_out <= 16'h8FE4	;
				14'b11010100100010: Data_out <= 16'h8FEA	;
				14'b11010100100011: Data_out <= 16'h8FF0	;
				14'b11010100100100: Data_out <= 16'h8FF6	;
				14'b11010100100101: Data_out <= 16'h8FFC	;
				14'b11010100100110: Data_out <= 16'h9002	;
				14'b11010100100111: Data_out <= 16'h9008	;
				14'b11010100101000: Data_out <= 16'h900F	;
				14'b11010100101001: Data_out <= 16'h9015	;
				14'b11010100101010: Data_out <= 16'h901B	;
				14'b11010100101011: Data_out <= 16'h9021	;
				14'b11010100101100: Data_out <= 16'h9027	;
				14'b11010100101101: Data_out <= 16'h902D	;
				14'b11010100101110: Data_out <= 16'h9033	;
				14'b11010100101111: Data_out <= 16'h9039	;
				14'b11010100110000: Data_out <= 16'h903F	;
				14'b11010100110001: Data_out <= 16'h9046	;
				14'b11010100110010: Data_out <= 16'h904C	;
				14'b11010100110011: Data_out <= 16'h9052	;
				14'b11010100110100: Data_out <= 16'h9058	;
				14'b11010100110101: Data_out <= 16'h905E	;
				14'b11010100110110: Data_out <= 16'h9064	;
				14'b11010100110111: Data_out <= 16'h906A	;
				14'b11010100111000: Data_out <= 16'h9071	;
				14'b11010100111001: Data_out <= 16'h9077	;
				14'b11010100111010: Data_out <= 16'h907D	;
				14'b11010100111011: Data_out <= 16'h9083	;
				14'b11010100111100: Data_out <= 16'h9089	;
				14'b11010100111101: Data_out <= 16'h908F	;
				14'b11010100111110: Data_out <= 16'h9096	;
				14'b11010100111111: Data_out <= 16'h909C	;
				14'b11010101000000: Data_out <= 16'h90A2	;
				14'b11010101000001: Data_out <= 16'h90A8	;
				14'b11010101000010: Data_out <= 16'h90AE	;
				14'b11010101000011: Data_out <= 16'h90B5	;
				14'b11010101000100: Data_out <= 16'h90BB	;
				14'b11010101000101: Data_out <= 16'h90C1	;
				14'b11010101000110: Data_out <= 16'h90C7	;
				14'b11010101000111: Data_out <= 16'h90CD	;
				14'b11010101001000: Data_out <= 16'h90D4	;
				14'b11010101001001: Data_out <= 16'h90DA	;
				14'b11010101001010: Data_out <= 16'h90E0	;
				14'b11010101001011: Data_out <= 16'h90E6	;
				14'b11010101001100: Data_out <= 16'h90ED	;
				14'b11010101001101: Data_out <= 16'h90F3	;
				14'b11010101001110: Data_out <= 16'h90F9	;
				14'b11010101001111: Data_out <= 16'h90FF	;
				14'b11010101010000: Data_out <= 16'h9106	;
				14'b11010101010001: Data_out <= 16'h910C	;
				14'b11010101010010: Data_out <= 16'h9112	;
				14'b11010101010011: Data_out <= 16'h9118	;
				14'b11010101010100: Data_out <= 16'h911F	;
				14'b11010101010101: Data_out <= 16'h9125	;
				14'b11010101010110: Data_out <= 16'h912B	;
				14'b11010101010111: Data_out <= 16'h9132	;
				14'b11010101011000: Data_out <= 16'h9138	;
				14'b11010101011001: Data_out <= 16'h913E	;
				14'b11010101011010: Data_out <= 16'h9144	;
				14'b11010101011011: Data_out <= 16'h914B	;
				14'b11010101011100: Data_out <= 16'h9151	;
				14'b11010101011101: Data_out <= 16'h9157	;
				14'b11010101011110: Data_out <= 16'h915E	;
				14'b11010101011111: Data_out <= 16'h9164	;
				14'b11010101100000: Data_out <= 16'h916A	;
				14'b11010101100001: Data_out <= 16'h9171	;
				14'b11010101100010: Data_out <= 16'h9177	;
				14'b11010101100011: Data_out <= 16'h917D	;
				14'b11010101100100: Data_out <= 16'h9184	;
				14'b11010101100101: Data_out <= 16'h918A	;
				14'b11010101100110: Data_out <= 16'h9190	;
				14'b11010101100111: Data_out <= 16'h9197	;
				14'b11010101101000: Data_out <= 16'h919D	;
				14'b11010101101001: Data_out <= 16'h91A3	;
				14'b11010101101010: Data_out <= 16'h91AA	;
				14'b11010101101011: Data_out <= 16'h91B0	;
				14'b11010101101100: Data_out <= 16'h91B7	;
				14'b11010101101101: Data_out <= 16'h91BD	;
				14'b11010101101110: Data_out <= 16'h91C3	;
				14'b11010101101111: Data_out <= 16'h91CA	;
				14'b11010101110000: Data_out <= 16'h91D0	;
				14'b11010101110001: Data_out <= 16'h91D6	;
				14'b11010101110010: Data_out <= 16'h91DD	;
				14'b11010101110011: Data_out <= 16'h91E3	;
				14'b11010101110100: Data_out <= 16'h91EA	;
				14'b11010101110101: Data_out <= 16'h91F0	;
				14'b11010101110110: Data_out <= 16'h91F7	;
				14'b11010101110111: Data_out <= 16'h91FD	;
				14'b11010101111000: Data_out <= 16'h9203	;
				14'b11010101111001: Data_out <= 16'h920A	;
				14'b11010101111010: Data_out <= 16'h9210	;
				14'b11010101111011: Data_out <= 16'h9217	;
				14'b11010101111100: Data_out <= 16'h921D	;
				14'b11010101111101: Data_out <= 16'h9224	;
				14'b11010101111110: Data_out <= 16'h922A	;
				14'b11010101111111: Data_out <= 16'h9230	;
				14'b11010110000000: Data_out <= 16'h9237	;
				14'b11010110000001: Data_out <= 16'h923D	;
				14'b11010110000010: Data_out <= 16'h9244	;
				14'b11010110000011: Data_out <= 16'h924A	;
				14'b11010110000100: Data_out <= 16'h9251	;
				14'b11010110000101: Data_out <= 16'h9257	;
				14'b11010110000110: Data_out <= 16'h925E	;
				14'b11010110000111: Data_out <= 16'h9264	;
				14'b11010110001000: Data_out <= 16'h926B	;
				14'b11010110001001: Data_out <= 16'h9271	;
				14'b11010110001010: Data_out <= 16'h9278	;
				14'b11010110001011: Data_out <= 16'h927E	;
				14'b11010110001100: Data_out <= 16'h9285	;
				14'b11010110001101: Data_out <= 16'h928B	;
				14'b11010110001110: Data_out <= 16'h9292	;
				14'b11010110001111: Data_out <= 16'h9298	;
				14'b11010110010000: Data_out <= 16'h929F	;
				14'b11010110010001: Data_out <= 16'h92A5	;
				14'b11010110010010: Data_out <= 16'h92AC	;
				14'b11010110010011: Data_out <= 16'h92B2	;
				14'b11010110010100: Data_out <= 16'h92B9	;
				14'b11010110010101: Data_out <= 16'h92BF	;
				14'b11010110010110: Data_out <= 16'h92C6	;
				14'b11010110010111: Data_out <= 16'h92CD	;
				14'b11010110011000: Data_out <= 16'h92D3	;
				14'b11010110011001: Data_out <= 16'h92DA	;
				14'b11010110011010: Data_out <= 16'h92E0	;
				14'b11010110011011: Data_out <= 16'h92E7	;
				14'b11010110011100: Data_out <= 16'h92ED	;
				14'b11010110011101: Data_out <= 16'h92F4	;
				14'b11010110011110: Data_out <= 16'h92FB	;
				14'b11010110011111: Data_out <= 16'h9301	;
				14'b11010110100000: Data_out <= 16'h9308	;
				14'b11010110100001: Data_out <= 16'h930E	;
				14'b11010110100010: Data_out <= 16'h9315	;
				14'b11010110100011: Data_out <= 16'h931C	;
				14'b11010110100100: Data_out <= 16'h9322	;
				14'b11010110100101: Data_out <= 16'h9329	;
				14'b11010110100110: Data_out <= 16'h932F	;
				14'b11010110100111: Data_out <= 16'h9336	;
				14'b11010110101000: Data_out <= 16'h933D	;
				14'b11010110101001: Data_out <= 16'h9343	;
				14'b11010110101010: Data_out <= 16'h934A	;
				14'b11010110101011: Data_out <= 16'h9351	;
				14'b11010110101100: Data_out <= 16'h9357	;
				14'b11010110101101: Data_out <= 16'h935E	;
				14'b11010110101110: Data_out <= 16'h9364	;
				14'b11010110101111: Data_out <= 16'h936B	;
				14'b11010110110000: Data_out <= 16'h9372	;
				14'b11010110110001: Data_out <= 16'h9378	;
				14'b11010110110010: Data_out <= 16'h937F	;
				14'b11010110110011: Data_out <= 16'h9386	;
				14'b11010110110100: Data_out <= 16'h938C	;
				14'b11010110110101: Data_out <= 16'h9393	;
				14'b11010110110110: Data_out <= 16'h939A	;
				14'b11010110110111: Data_out <= 16'h93A0	;
				14'b11010110111000: Data_out <= 16'h93A7	;
				14'b11010110111001: Data_out <= 16'h93AE	;
				14'b11010110111010: Data_out <= 16'h93B5	;
				14'b11010110111011: Data_out <= 16'h93BB	;
				14'b11010110111100: Data_out <= 16'h93C2	;
				14'b11010110111101: Data_out <= 16'h93C9	;
				14'b11010110111110: Data_out <= 16'h93CF	;
				14'b11010110111111: Data_out <= 16'h93D6	;
				14'b11010111000000: Data_out <= 16'h93DD	;
				14'b11010111000001: Data_out <= 16'h93E4	;
				14'b11010111000010: Data_out <= 16'h93EA	;
				14'b11010111000011: Data_out <= 16'h93F1	;
				14'b11010111000100: Data_out <= 16'h93F8	;
				14'b11010111000101: Data_out <= 16'h93FE	;
				14'b11010111000110: Data_out <= 16'h9405	;
				14'b11010111000111: Data_out <= 16'h940C	;
				14'b11010111001000: Data_out <= 16'h9413	;
				14'b11010111001001: Data_out <= 16'h9419	;
				14'b11010111001010: Data_out <= 16'h9420	;
				14'b11010111001011: Data_out <= 16'h9427	;
				14'b11010111001100: Data_out <= 16'h942E	;
				14'b11010111001101: Data_out <= 16'h9435	;
				14'b11010111001110: Data_out <= 16'h943B	;
				14'b11010111001111: Data_out <= 16'h9442	;
				14'b11010111010000: Data_out <= 16'h9449	;
				14'b11010111010001: Data_out <= 16'h9450	;
				14'b11010111010010: Data_out <= 16'h9456	;
				14'b11010111010011: Data_out <= 16'h945D	;
				14'b11010111010100: Data_out <= 16'h9464	;
				14'b11010111010101: Data_out <= 16'h946B	;
				14'b11010111010110: Data_out <= 16'h9472	;
				14'b11010111010111: Data_out <= 16'h9478	;
				14'b11010111011000: Data_out <= 16'h947F	;
				14'b11010111011001: Data_out <= 16'h9486	;
				14'b11010111011010: Data_out <= 16'h948D	;
				14'b11010111011011: Data_out <= 16'h9494	;
				14'b11010111011100: Data_out <= 16'h949B	;
				14'b11010111011101: Data_out <= 16'h94A1	;
				14'b11010111011110: Data_out <= 16'h94A8	;
				14'b11010111011111: Data_out <= 16'h94AF	;
				14'b11010111100000: Data_out <= 16'h94B6	;
				14'b11010111100001: Data_out <= 16'h94BD	;
				14'b11010111100010: Data_out <= 16'h94C4	;
				14'b11010111100011: Data_out <= 16'h94CB	;
				14'b11010111100100: Data_out <= 16'h94D1	;
				14'b11010111100101: Data_out <= 16'h94D8	;
				14'b11010111100110: Data_out <= 16'h94DF	;
				14'b11010111100111: Data_out <= 16'h94E6	;
				14'b11010111101000: Data_out <= 16'h94ED	;
				14'b11010111101001: Data_out <= 16'h94F4	;
				14'b11010111101010: Data_out <= 16'h94FB	;
				14'b11010111101011: Data_out <= 16'h9502	;
				14'b11010111101100: Data_out <= 16'h9509	;
				14'b11010111101101: Data_out <= 16'h950F	;
				14'b11010111101110: Data_out <= 16'h9516	;
				14'b11010111101111: Data_out <= 16'h951D	;
				14'b11010111110000: Data_out <= 16'h9524	;
				14'b11010111110001: Data_out <= 16'h952B	;
				14'b11010111110010: Data_out <= 16'h9532	;
				14'b11010111110011: Data_out <= 16'h9539	;
				14'b11010111110100: Data_out <= 16'h9540	;
				14'b11010111110101: Data_out <= 16'h9547	;
				14'b11010111110110: Data_out <= 16'h954E	;
				14'b11010111110111: Data_out <= 16'h9555	;
				14'b11010111111000: Data_out <= 16'h955C	;
				14'b11010111111001: Data_out <= 16'h9563	;
				14'b11010111111010: Data_out <= 16'h956A	;
				14'b11010111111011: Data_out <= 16'h9570	;
				14'b11010111111100: Data_out <= 16'h9577	;
				14'b11010111111101: Data_out <= 16'h957E	;
				14'b11010111111110: Data_out <= 16'h9585	;
				14'b11010111111111: Data_out <= 16'h958C	;
				14'b11011000000000: Data_out <= 16'h9593	;
				14'b11011000000001: Data_out <= 16'h959A	;
				14'b11011000000010: Data_out <= 16'h95A1	;
				14'b11011000000011: Data_out <= 16'h95A8	;
				14'b11011000000100: Data_out <= 16'h95AF	;
				14'b11011000000101: Data_out <= 16'h95B6	;
				14'b11011000000110: Data_out <= 16'h95BD	;
				14'b11011000000111: Data_out <= 16'h95C4	;
				14'b11011000001000: Data_out <= 16'h95CB	;
				14'b11011000001001: Data_out <= 16'h95D2	;
				14'b11011000001010: Data_out <= 16'h95D9	;
				14'b11011000001011: Data_out <= 16'h95E0	;
				14'b11011000001100: Data_out <= 16'h95E7	;
				14'b11011000001101: Data_out <= 16'h95EE	;
				14'b11011000001110: Data_out <= 16'h95F5	;
				14'b11011000001111: Data_out <= 16'h95FD	;
				14'b11011000010000: Data_out <= 16'h9604	;
				14'b11011000010001: Data_out <= 16'h960B	;
				14'b11011000010010: Data_out <= 16'h9612	;
				14'b11011000010011: Data_out <= 16'h9619	;
				14'b11011000010100: Data_out <= 16'h9620	;
				14'b11011000010101: Data_out <= 16'h9627	;
				14'b11011000010110: Data_out <= 16'h962E	;
				14'b11011000010111: Data_out <= 16'h9635	;
				14'b11011000011000: Data_out <= 16'h963C	;
				14'b11011000011001: Data_out <= 16'h9643	;
				14'b11011000011010: Data_out <= 16'h964A	;
				14'b11011000011011: Data_out <= 16'h9651	;
				14'b11011000011100: Data_out <= 16'h9658	;
				14'b11011000011101: Data_out <= 16'h965F	;
				14'b11011000011110: Data_out <= 16'h9667	;
				14'b11011000011111: Data_out <= 16'h966E	;
				14'b11011000100000: Data_out <= 16'h9675	;
				14'b11011000100001: Data_out <= 16'h967C	;
				14'b11011000100010: Data_out <= 16'h9683	;
				14'b11011000100011: Data_out <= 16'h968A	;
				14'b11011000100100: Data_out <= 16'h9691	;
				14'b11011000100101: Data_out <= 16'h9698	;
				14'b11011000100110: Data_out <= 16'h96A0	;
				14'b11011000100111: Data_out <= 16'h96A7	;
				14'b11011000101000: Data_out <= 16'h96AE	;
				14'b11011000101001: Data_out <= 16'h96B5	;
				14'b11011000101010: Data_out <= 16'h96BC	;
				14'b11011000101011: Data_out <= 16'h96C3	;
				14'b11011000101100: Data_out <= 16'h96CA	;
				14'b11011000101101: Data_out <= 16'h96D2	;
				14'b11011000101110: Data_out <= 16'h96D9	;
				14'b11011000101111: Data_out <= 16'h96E0	;
				14'b11011000110000: Data_out <= 16'h96E7	;
				14'b11011000110001: Data_out <= 16'h96EE	;
				14'b11011000110010: Data_out <= 16'h96F5	;
				14'b11011000110011: Data_out <= 16'h96FD	;
				14'b11011000110100: Data_out <= 16'h9704	;
				14'b11011000110101: Data_out <= 16'h970B	;
				14'b11011000110110: Data_out <= 16'h9712	;
				14'b11011000110111: Data_out <= 16'h9719	;
				14'b11011000111000: Data_out <= 16'h9721	;
				14'b11011000111001: Data_out <= 16'h9728	;
				14'b11011000111010: Data_out <= 16'h972F	;
				14'b11011000111011: Data_out <= 16'h9736	;
				14'b11011000111100: Data_out <= 16'h973D	;
				14'b11011000111101: Data_out <= 16'h9745	;
				14'b11011000111110: Data_out <= 16'h974C	;
				14'b11011000111111: Data_out <= 16'h9753	;
				14'b11011001000000: Data_out <= 16'h975A	;
				14'b11011001000001: Data_out <= 16'h9762	;
				14'b11011001000010: Data_out <= 16'h9769	;
				14'b11011001000011: Data_out <= 16'h9770	;
				14'b11011001000100: Data_out <= 16'h9777	;
				14'b11011001000101: Data_out <= 16'h977F	;
				14'b11011001000110: Data_out <= 16'h9786	;
				14'b11011001000111: Data_out <= 16'h978D	;
				14'b11011001001000: Data_out <= 16'h9794	;
				14'b11011001001001: Data_out <= 16'h979C	;
				14'b11011001001010: Data_out <= 16'h97A3	;
				14'b11011001001011: Data_out <= 16'h97AA	;
				14'b11011001001100: Data_out <= 16'h97B1	;
				14'b11011001001101: Data_out <= 16'h97B9	;
				14'b11011001001110: Data_out <= 16'h97C0	;
				14'b11011001001111: Data_out <= 16'h97C7	;
				14'b11011001010000: Data_out <= 16'h97CF	;
				14'b11011001010001: Data_out <= 16'h97D6	;
				14'b11011001010010: Data_out <= 16'h97DD	;
				14'b11011001010011: Data_out <= 16'h97E4	;
				14'b11011001010100: Data_out <= 16'h97EC	;
				14'b11011001010101: Data_out <= 16'h97F3	;
				14'b11011001010110: Data_out <= 16'h97FA	;
				14'b11011001010111: Data_out <= 16'h9802	;
				14'b11011001011000: Data_out <= 16'h9809	;
				14'b11011001011001: Data_out <= 16'h9810	;
				14'b11011001011010: Data_out <= 16'h9818	;
				14'b11011001011011: Data_out <= 16'h981F	;
				14'b11011001011100: Data_out <= 16'h9826	;
				14'b11011001011101: Data_out <= 16'h982E	;
				14'b11011001011110: Data_out <= 16'h9835	;
				14'b11011001011111: Data_out <= 16'h983C	;
				14'b11011001100000: Data_out <= 16'h9844	;
				14'b11011001100001: Data_out <= 16'h984B	;
				14'b11011001100010: Data_out <= 16'h9853	;
				14'b11011001100011: Data_out <= 16'h985A	;
				14'b11011001100100: Data_out <= 16'h9861	;
				14'b11011001100101: Data_out <= 16'h9869	;
				14'b11011001100110: Data_out <= 16'h9870	;
				14'b11011001100111: Data_out <= 16'h9877	;
				14'b11011001101000: Data_out <= 16'h987F	;
				14'b11011001101001: Data_out <= 16'h9886	;
				14'b11011001101010: Data_out <= 16'h988E	;
				14'b11011001101011: Data_out <= 16'h9895	;
				14'b11011001101100: Data_out <= 16'h989C	;
				14'b11011001101101: Data_out <= 16'h98A4	;
				14'b11011001101110: Data_out <= 16'h98AB	;
				14'b11011001101111: Data_out <= 16'h98B3	;
				14'b11011001110000: Data_out <= 16'h98BA	;
				14'b11011001110001: Data_out <= 16'h98C2	;
				14'b11011001110010: Data_out <= 16'h98C9	;
				14'b11011001110011: Data_out <= 16'h98D0	;
				14'b11011001110100: Data_out <= 16'h98D8	;
				14'b11011001110101: Data_out <= 16'h98DF	;
				14'b11011001110110: Data_out <= 16'h98E7	;
				14'b11011001110111: Data_out <= 16'h98EE	;
				14'b11011001111000: Data_out <= 16'h98F6	;
				14'b11011001111001: Data_out <= 16'h98FD	;
				14'b11011001111010: Data_out <= 16'h9905	;
				14'b11011001111011: Data_out <= 16'h990C	;
				14'b11011001111100: Data_out <= 16'h9913	;
				14'b11011001111101: Data_out <= 16'h991B	;
				14'b11011001111110: Data_out <= 16'h9922	;
				14'b11011001111111: Data_out <= 16'h992A	;
				14'b11011010000000: Data_out <= 16'h9931	;
				14'b11011010000001: Data_out <= 16'h9939	;
				14'b11011010000010: Data_out <= 16'h9940	;
				14'b11011010000011: Data_out <= 16'h9948	;
				14'b11011010000100: Data_out <= 16'h994F	;
				14'b11011010000101: Data_out <= 16'h9957	;
				14'b11011010000110: Data_out <= 16'h995E	;
				14'b11011010000111: Data_out <= 16'h9966	;
				14'b11011010001000: Data_out <= 16'h996D	;
				14'b11011010001001: Data_out <= 16'h9975	;
				14'b11011010001010: Data_out <= 16'h997C	;
				14'b11011010001011: Data_out <= 16'h9984	;
				14'b11011010001100: Data_out <= 16'h998C	;
				14'b11011010001101: Data_out <= 16'h9993	;
				14'b11011010001110: Data_out <= 16'h999B	;
				14'b11011010001111: Data_out <= 16'h99A2	;
				14'b11011010010000: Data_out <= 16'h99AA	;
				14'b11011010010001: Data_out <= 16'h99B1	;
				14'b11011010010010: Data_out <= 16'h99B9	;
				14'b11011010010011: Data_out <= 16'h99C0	;
				14'b11011010010100: Data_out <= 16'h99C8	;
				14'b11011010010101: Data_out <= 16'h99CF	;
				14'b11011010010110: Data_out <= 16'h99D7	;
				14'b11011010010111: Data_out <= 16'h99DF	;
				14'b11011010011000: Data_out <= 16'h99E6	;
				14'b11011010011001: Data_out <= 16'h99EE	;
				14'b11011010011010: Data_out <= 16'h99F5	;
				14'b11011010011011: Data_out <= 16'h99FD	;
				14'b11011010011100: Data_out <= 16'h9A05	;
				14'b11011010011101: Data_out <= 16'h9A0C	;
				14'b11011010011110: Data_out <= 16'h9A14	;
				14'b11011010011111: Data_out <= 16'h9A1B	;
				14'b11011010100000: Data_out <= 16'h9A23	;
				14'b11011010100001: Data_out <= 16'h9A2B	;
				14'b11011010100010: Data_out <= 16'h9A32	;
				14'b11011010100011: Data_out <= 16'h9A3A	;
				14'b11011010100100: Data_out <= 16'h9A41	;
				14'b11011010100101: Data_out <= 16'h9A49	;
				14'b11011010100110: Data_out <= 16'h9A51	;
				14'b11011010100111: Data_out <= 16'h9A58	;
				14'b11011010101000: Data_out <= 16'h9A60	;
				14'b11011010101001: Data_out <= 16'h9A68	;
				14'b11011010101010: Data_out <= 16'h9A6F	;
				14'b11011010101011: Data_out <= 16'h9A77	;
				14'b11011010101100: Data_out <= 16'h9A7E	;
				14'b11011010101101: Data_out <= 16'h9A86	;
				14'b11011010101110: Data_out <= 16'h9A8E	;
				14'b11011010101111: Data_out <= 16'h9A95	;
				14'b11011010110000: Data_out <= 16'h9A9D	;
				14'b11011010110001: Data_out <= 16'h9AA5	;
				14'b11011010110010: Data_out <= 16'h9AAC	;
				14'b11011010110011: Data_out <= 16'h9AB4	;
				14'b11011010110100: Data_out <= 16'h9ABC	;
				14'b11011010110101: Data_out <= 16'h9AC4	;
				14'b11011010110110: Data_out <= 16'h9ACB	;
				14'b11011010110111: Data_out <= 16'h9AD3	;
				14'b11011010111000: Data_out <= 16'h9ADB	;
				14'b11011010111001: Data_out <= 16'h9AE2	;
				14'b11011010111010: Data_out <= 16'h9AEA	;
				14'b11011010111011: Data_out <= 16'h9AF2	;
				14'b11011010111100: Data_out <= 16'h9AF9	;
				14'b11011010111101: Data_out <= 16'h9B01	;
				14'b11011010111110: Data_out <= 16'h9B09	;
				14'b11011010111111: Data_out <= 16'h9B11	;
				14'b11011011000000: Data_out <= 16'h9B18	;
				14'b11011011000001: Data_out <= 16'h9B20	;
				14'b11011011000010: Data_out <= 16'h9B28	;
				14'b11011011000011: Data_out <= 16'h9B30	;
				14'b11011011000100: Data_out <= 16'h9B37	;
				14'b11011011000101: Data_out <= 16'h9B3F	;
				14'b11011011000110: Data_out <= 16'h9B47	;
				14'b11011011000111: Data_out <= 16'h9B4F	;
				14'b11011011001000: Data_out <= 16'h9B56	;
				14'b11011011001001: Data_out <= 16'h9B5E	;
				14'b11011011001010: Data_out <= 16'h9B66	;
				14'b11011011001011: Data_out <= 16'h9B6E	;
				14'b11011011001100: Data_out <= 16'h9B75	;
				14'b11011011001101: Data_out <= 16'h9B7D	;
				14'b11011011001110: Data_out <= 16'h9B85	;
				14'b11011011001111: Data_out <= 16'h9B8D	;
				14'b11011011010000: Data_out <= 16'h9B95	;
				14'b11011011010001: Data_out <= 16'h9B9C	;
				14'b11011011010010: Data_out <= 16'h9BA4	;
				14'b11011011010011: Data_out <= 16'h9BAC	;
				14'b11011011010100: Data_out <= 16'h9BB4	;
				14'b11011011010101: Data_out <= 16'h9BBC	;
				14'b11011011010110: Data_out <= 16'h9BC3	;
				14'b11011011010111: Data_out <= 16'h9BCB	;
				14'b11011011011000: Data_out <= 16'h9BD3	;
				14'b11011011011001: Data_out <= 16'h9BDB	;
				14'b11011011011010: Data_out <= 16'h9BE3	;
				14'b11011011011011: Data_out <= 16'h9BEA	;
				14'b11011011011100: Data_out <= 16'h9BF2	;
				14'b11011011011101: Data_out <= 16'h9BFA	;
				14'b11011011011110: Data_out <= 16'h9C02	;
				14'b11011011011111: Data_out <= 16'h9C0A	;
				14'b11011011100000: Data_out <= 16'h9C12	;
				14'b11011011100001: Data_out <= 16'h9C1A	;
				14'b11011011100010: Data_out <= 16'h9C21	;
				14'b11011011100011: Data_out <= 16'h9C29	;
				14'b11011011100100: Data_out <= 16'h9C31	;
				14'b11011011100101: Data_out <= 16'h9C39	;
				14'b11011011100110: Data_out <= 16'h9C41	;
				14'b11011011100111: Data_out <= 16'h9C49	;
				14'b11011011101000: Data_out <= 16'h9C51	;
				14'b11011011101001: Data_out <= 16'h9C59	;
				14'b11011011101010: Data_out <= 16'h9C60	;
				14'b11011011101011: Data_out <= 16'h9C68	;
				14'b11011011101100: Data_out <= 16'h9C70	;
				14'b11011011101101: Data_out <= 16'h9C78	;
				14'b11011011101110: Data_out <= 16'h9C80	;
				14'b11011011101111: Data_out <= 16'h9C88	;
				14'b11011011110000: Data_out <= 16'h9C90	;
				14'b11011011110001: Data_out <= 16'h9C98	;
				14'b11011011110010: Data_out <= 16'h9CA0	;
				14'b11011011110011: Data_out <= 16'h9CA8	;
				14'b11011011110100: Data_out <= 16'h9CAF	;
				14'b11011011110101: Data_out <= 16'h9CB7	;
				14'b11011011110110: Data_out <= 16'h9CBF	;
				14'b11011011110111: Data_out <= 16'h9CC7	;
				14'b11011011111000: Data_out <= 16'h9CCF	;
				14'b11011011111001: Data_out <= 16'h9CD7	;
				14'b11011011111010: Data_out <= 16'h9CDF	;
				14'b11011011111011: Data_out <= 16'h9CE7	;
				14'b11011011111100: Data_out <= 16'h9CEF	;
				14'b11011011111101: Data_out <= 16'h9CF7	;
				14'b11011011111110: Data_out <= 16'h9CFF	;
				14'b11011011111111: Data_out <= 16'h9D07	;
				14'b11011100000000: Data_out <= 16'h9D0F	;
				14'b11011100000001: Data_out <= 16'h9D17	;
				14'b11011100000010: Data_out <= 16'h9D1F	;
				14'b11011100000011: Data_out <= 16'h9D27	;
				14'b11011100000100: Data_out <= 16'h9D2F	;
				14'b11011100000101: Data_out <= 16'h9D37	;
				14'b11011100000110: Data_out <= 16'h9D3F	;
				14'b11011100000111: Data_out <= 16'h9D47	;
				14'b11011100001000: Data_out <= 16'h9D4F	;
				14'b11011100001001: Data_out <= 16'h9D57	;
				14'b11011100001010: Data_out <= 16'h9D5F	;
				14'b11011100001011: Data_out <= 16'h9D67	;
				14'b11011100001100: Data_out <= 16'h9D6F	;
				14'b11011100001101: Data_out <= 16'h9D77	;
				14'b11011100001110: Data_out <= 16'h9D7F	;
				14'b11011100001111: Data_out <= 16'h9D87	;
				14'b11011100010000: Data_out <= 16'h9D8F	;
				14'b11011100010001: Data_out <= 16'h9D97	;
				14'b11011100010010: Data_out <= 16'h9D9F	;
				14'b11011100010011: Data_out <= 16'h9DA7	;
				14'b11011100010100: Data_out <= 16'h9DAF	;
				14'b11011100010101: Data_out <= 16'h9DB7	;
				14'b11011100010110: Data_out <= 16'h9DBF	;
				14'b11011100010111: Data_out <= 16'h9DC7	;
				14'b11011100011000: Data_out <= 16'h9DCF	;
				14'b11011100011001: Data_out <= 16'h9DD7	;
				14'b11011100011010: Data_out <= 16'h9DDF	;
				14'b11011100011011: Data_out <= 16'h9DE7	;
				14'b11011100011100: Data_out <= 16'h9DF0	;
				14'b11011100011101: Data_out <= 16'h9DF8	;
				14'b11011100011110: Data_out <= 16'h9E00	;
				14'b11011100011111: Data_out <= 16'h9E08	;
				14'b11011100100000: Data_out <= 16'h9E10	;
				14'b11011100100001: Data_out <= 16'h9E18	;
				14'b11011100100010: Data_out <= 16'h9E20	;
				14'b11011100100011: Data_out <= 16'h9E28	;
				14'b11011100100100: Data_out <= 16'h9E30	;
				14'b11011100100101: Data_out <= 16'h9E38	;
				14'b11011100100110: Data_out <= 16'h9E40	;
				14'b11011100100111: Data_out <= 16'h9E49	;
				14'b11011100101000: Data_out <= 16'h9E51	;
				14'b11011100101001: Data_out <= 16'h9E59	;
				14'b11011100101010: Data_out <= 16'h9E61	;
				14'b11011100101011: Data_out <= 16'h9E69	;
				14'b11011100101100: Data_out <= 16'h9E71	;
				14'b11011100101101: Data_out <= 16'h9E79	;
				14'b11011100101110: Data_out <= 16'h9E81	;
				14'b11011100101111: Data_out <= 16'h9E8A	;
				14'b11011100110000: Data_out <= 16'h9E92	;
				14'b11011100110001: Data_out <= 16'h9E9A	;
				14'b11011100110010: Data_out <= 16'h9EA2	;
				14'b11011100110011: Data_out <= 16'h9EAA	;
				14'b11011100110100: Data_out <= 16'h9EB2	;
				14'b11011100110101: Data_out <= 16'h9EBB	;
				14'b11011100110110: Data_out <= 16'h9EC3	;
				14'b11011100110111: Data_out <= 16'h9ECB	;
				14'b11011100111000: Data_out <= 16'h9ED3	;
				14'b11011100111001: Data_out <= 16'h9EDB	;
				14'b11011100111010: Data_out <= 16'h9EE3	;
				14'b11011100111011: Data_out <= 16'h9EEC	;
				14'b11011100111100: Data_out <= 16'h9EF4	;
				14'b11011100111101: Data_out <= 16'h9EFC	;
				14'b11011100111110: Data_out <= 16'h9F04	;
				14'b11011100111111: Data_out <= 16'h9F0C	;
				14'b11011101000000: Data_out <= 16'h9F15	;
				14'b11011101000001: Data_out <= 16'h9F1D	;
				14'b11011101000010: Data_out <= 16'h9F25	;
				14'b11011101000011: Data_out <= 16'h9F2D	;
				14'b11011101000100: Data_out <= 16'h9F35	;
				14'b11011101000101: Data_out <= 16'h9F3E	;
				14'b11011101000110: Data_out <= 16'h9F46	;
				14'b11011101000111: Data_out <= 16'h9F4E	;
				14'b11011101001000: Data_out <= 16'h9F56	;
				14'b11011101001001: Data_out <= 16'h9F5F	;
				14'b11011101001010: Data_out <= 16'h9F67	;
				14'b11011101001011: Data_out <= 16'h9F6F	;
				14'b11011101001100: Data_out <= 16'h9F77	;
				14'b11011101001101: Data_out <= 16'h9F80	;
				14'b11011101001110: Data_out <= 16'h9F88	;
				14'b11011101001111: Data_out <= 16'h9F90	;
				14'b11011101010000: Data_out <= 16'h9F98	;
				14'b11011101010001: Data_out <= 16'h9FA1	;
				14'b11011101010010: Data_out <= 16'h9FA9	;
				14'b11011101010011: Data_out <= 16'h9FB1	;
				14'b11011101010100: Data_out <= 16'h9FBA	;
				14'b11011101010101: Data_out <= 16'h9FC2	;
				14'b11011101010110: Data_out <= 16'h9FCA	;
				14'b11011101010111: Data_out <= 16'h9FD2	;
				14'b11011101011000: Data_out <= 16'h9FDB	;
				14'b11011101011001: Data_out <= 16'h9FE3	;
				14'b11011101011010: Data_out <= 16'h9FEB	;
				14'b11011101011011: Data_out <= 16'h9FF4	;
				14'b11011101011100: Data_out <= 16'h9FFC	;
				14'b11011101011101: Data_out <= 16'hA004	;
				14'b11011101011110: Data_out <= 16'hA00D	;
				14'b11011101011111: Data_out <= 16'hA015	;
				14'b11011101100000: Data_out <= 16'hA01D	;
				14'b11011101100001: Data_out <= 16'hA025	;
				14'b11011101100010: Data_out <= 16'hA02E	;
				14'b11011101100011: Data_out <= 16'hA036	;
				14'b11011101100100: Data_out <= 16'hA03E	;
				14'b11011101100101: Data_out <= 16'hA047	;
				14'b11011101100110: Data_out <= 16'hA04F	;
				14'b11011101100111: Data_out <= 16'hA058	;
				14'b11011101101000: Data_out <= 16'hA060	;
				14'b11011101101001: Data_out <= 16'hA068	;
				14'b11011101101010: Data_out <= 16'hA071	;
				14'b11011101101011: Data_out <= 16'hA079	;
				14'b11011101101100: Data_out <= 16'hA081	;
				14'b11011101101101: Data_out <= 16'hA08A	;
				14'b11011101101110: Data_out <= 16'hA092	;
				14'b11011101101111: Data_out <= 16'hA09A	;
				14'b11011101110000: Data_out <= 16'hA0A3	;
				14'b11011101110001: Data_out <= 16'hA0AB	;
				14'b11011101110010: Data_out <= 16'hA0B4	;
				14'b11011101110011: Data_out <= 16'hA0BC	;
				14'b11011101110100: Data_out <= 16'hA0C4	;
				14'b11011101110101: Data_out <= 16'hA0CD	;
				14'b11011101110110: Data_out <= 16'hA0D5	;
				14'b11011101110111: Data_out <= 16'hA0DE	;
				14'b11011101111000: Data_out <= 16'hA0E6	;
				14'b11011101111001: Data_out <= 16'hA0EE	;
				14'b11011101111010: Data_out <= 16'hA0F7	;
				14'b11011101111011: Data_out <= 16'hA0FF	;
				14'b11011101111100: Data_out <= 16'hA108	;
				14'b11011101111101: Data_out <= 16'hA110	;
				14'b11011101111110: Data_out <= 16'hA118	;
				14'b11011101111111: Data_out <= 16'hA121	;
				14'b11011110000000: Data_out <= 16'hA129	;
				14'b11011110000001: Data_out <= 16'hA132	;
				14'b11011110000010: Data_out <= 16'hA13A	;
				14'b11011110000011: Data_out <= 16'hA143	;
				14'b11011110000100: Data_out <= 16'hA14B	;
				14'b11011110000101: Data_out <= 16'hA154	;
				14'b11011110000110: Data_out <= 16'hA15C	;
				14'b11011110000111: Data_out <= 16'hA165	;
				14'b11011110001000: Data_out <= 16'hA16D	;
				14'b11011110001001: Data_out <= 16'hA175	;
				14'b11011110001010: Data_out <= 16'hA17E	;
				14'b11011110001011: Data_out <= 16'hA186	;
				14'b11011110001100: Data_out <= 16'hA18F	;
				14'b11011110001101: Data_out <= 16'hA197	;
				14'b11011110001110: Data_out <= 16'hA1A0	;
				14'b11011110001111: Data_out <= 16'hA1A8	;
				14'b11011110010000: Data_out <= 16'hA1B1	;
				14'b11011110010001: Data_out <= 16'hA1B9	;
				14'b11011110010010: Data_out <= 16'hA1C2	;
				14'b11011110010011: Data_out <= 16'hA1CA	;
				14'b11011110010100: Data_out <= 16'hA1D3	;
				14'b11011110010101: Data_out <= 16'hA1DB	;
				14'b11011110010110: Data_out <= 16'hA1E4	;
				14'b11011110010111: Data_out <= 16'hA1EC	;
				14'b11011110011000: Data_out <= 16'hA1F5	;
				14'b11011110011001: Data_out <= 16'hA1FD	;
				14'b11011110011010: Data_out <= 16'hA206	;
				14'b11011110011011: Data_out <= 16'hA20E	;
				14'b11011110011100: Data_out <= 16'hA217	;
				14'b11011110011101: Data_out <= 16'hA220	;
				14'b11011110011110: Data_out <= 16'hA228	;
				14'b11011110011111: Data_out <= 16'hA231	;
				14'b11011110100000: Data_out <= 16'hA239	;
				14'b11011110100001: Data_out <= 16'hA242	;
				14'b11011110100010: Data_out <= 16'hA24A	;
				14'b11011110100011: Data_out <= 16'hA253	;
				14'b11011110100100: Data_out <= 16'hA25B	;
				14'b11011110100101: Data_out <= 16'hA264	;
				14'b11011110100110: Data_out <= 16'hA26D	;
				14'b11011110100111: Data_out <= 16'hA275	;
				14'b11011110101000: Data_out <= 16'hA27E	;
				14'b11011110101001: Data_out <= 16'hA286	;
				14'b11011110101010: Data_out <= 16'hA28F	;
				14'b11011110101011: Data_out <= 16'hA298	;
				14'b11011110101100: Data_out <= 16'hA2A0	;
				14'b11011110101101: Data_out <= 16'hA2A9	;
				14'b11011110101110: Data_out <= 16'hA2B1	;
				14'b11011110101111: Data_out <= 16'hA2BA	;
				14'b11011110110000: Data_out <= 16'hA2C3	;
				14'b11011110110001: Data_out <= 16'hA2CB	;
				14'b11011110110010: Data_out <= 16'hA2D4	;
				14'b11011110110011: Data_out <= 16'hA2DC	;
				14'b11011110110100: Data_out <= 16'hA2E5	;
				14'b11011110110101: Data_out <= 16'hA2EE	;
				14'b11011110110110: Data_out <= 16'hA2F6	;
				14'b11011110110111: Data_out <= 16'hA2FF	;
				14'b11011110111000: Data_out <= 16'hA307	;
				14'b11011110111001: Data_out <= 16'hA310	;
				14'b11011110111010: Data_out <= 16'hA319	;
				14'b11011110111011: Data_out <= 16'hA321	;
				14'b11011110111100: Data_out <= 16'hA32A	;
				14'b11011110111101: Data_out <= 16'hA333	;
				14'b11011110111110: Data_out <= 16'hA33B	;
				14'b11011110111111: Data_out <= 16'hA344	;
				14'b11011111000000: Data_out <= 16'hA34D	;
				14'b11011111000001: Data_out <= 16'hA355	;
				14'b11011111000010: Data_out <= 16'hA35E	;
				14'b11011111000011: Data_out <= 16'hA367	;
				14'b11011111000100: Data_out <= 16'hA36F	;
				14'b11011111000101: Data_out <= 16'hA378	;
				14'b11011111000110: Data_out <= 16'hA381	;
				14'b11011111000111: Data_out <= 16'hA389	;
				14'b11011111001000: Data_out <= 16'hA392	;
				14'b11011111001001: Data_out <= 16'hA39B	;
				14'b11011111001010: Data_out <= 16'hA3A4	;
				14'b11011111001011: Data_out <= 16'hA3AC	;
				14'b11011111001100: Data_out <= 16'hA3B5	;
				14'b11011111001101: Data_out <= 16'hA3BE	;
				14'b11011111001110: Data_out <= 16'hA3C6	;
				14'b11011111001111: Data_out <= 16'hA3CF	;
				14'b11011111010000: Data_out <= 16'hA3D8	;
				14'b11011111010001: Data_out <= 16'hA3E0	;
				14'b11011111010010: Data_out <= 16'hA3E9	;
				14'b11011111010011: Data_out <= 16'hA3F2	;
				14'b11011111010100: Data_out <= 16'hA3FB	;
				14'b11011111010101: Data_out <= 16'hA403	;
				14'b11011111010110: Data_out <= 16'hA40C	;
				14'b11011111010111: Data_out <= 16'hA415	;
				14'b11011111011000: Data_out <= 16'hA41E	;
				14'b11011111011001: Data_out <= 16'hA426	;
				14'b11011111011010: Data_out <= 16'hA42F	;
				14'b11011111011011: Data_out <= 16'hA438	;
				14'b11011111011100: Data_out <= 16'hA441	;
				14'b11011111011101: Data_out <= 16'hA449	;
				14'b11011111011110: Data_out <= 16'hA452	;
				14'b11011111011111: Data_out <= 16'hA45B	;
				14'b11011111100000: Data_out <= 16'hA464	;
				14'b11011111100001: Data_out <= 16'hA46D	;
				14'b11011111100010: Data_out <= 16'hA475	;
				14'b11011111100011: Data_out <= 16'hA47E	;
				14'b11011111100100: Data_out <= 16'hA487	;
				14'b11011111100101: Data_out <= 16'hA490	;
				14'b11011111100110: Data_out <= 16'hA498	;
				14'b11011111100111: Data_out <= 16'hA4A1	;
				14'b11011111101000: Data_out <= 16'hA4AA	;
				14'b11011111101001: Data_out <= 16'hA4B3	;
				14'b11011111101010: Data_out <= 16'hA4BC	;
				14'b11011111101011: Data_out <= 16'hA4C4	;
				14'b11011111101100: Data_out <= 16'hA4CD	;
				14'b11011111101101: Data_out <= 16'hA4D6	;
				14'b11011111101110: Data_out <= 16'hA4DF	;
				14'b11011111101111: Data_out <= 16'hA4E8	;
				14'b11011111110000: Data_out <= 16'hA4F1	;
				14'b11011111110001: Data_out <= 16'hA4F9	;
				14'b11011111110010: Data_out <= 16'hA502	;
				14'b11011111110011: Data_out <= 16'hA50B	;
				14'b11011111110100: Data_out <= 16'hA514	;
				14'b11011111110101: Data_out <= 16'hA51D	;
				14'b11011111110110: Data_out <= 16'hA526	;
				14'b11011111110111: Data_out <= 16'hA52F	;
				14'b11011111111000: Data_out <= 16'hA537	;
				14'b11011111111001: Data_out <= 16'hA540	;
				14'b11011111111010: Data_out <= 16'hA549	;
				14'b11011111111011: Data_out <= 16'hA552	;
				14'b11011111111100: Data_out <= 16'hA55B	;
				14'b11011111111101: Data_out <= 16'hA564	;
				14'b11011111111110: Data_out <= 16'hA56D	;
				14'b11011111111111: Data_out <= 16'hA575	;
				14'b11100000000000: Data_out <= 16'hA57E	;
				14'b11100000000001: Data_out <= 16'hA587	;
				14'b11100000000010: Data_out <= 16'hA590	;
				14'b11100000000011: Data_out <= 16'hA599	;
				14'b11100000000100: Data_out <= 16'hA5A2	;
				14'b11100000000101: Data_out <= 16'hA5AB	;
				14'b11100000000110: Data_out <= 16'hA5B4	;
				14'b11100000000111: Data_out <= 16'hA5BD	;
				14'b11100000001000: Data_out <= 16'hA5C6	;
				14'b11100000001001: Data_out <= 16'hA5CE	;
				14'b11100000001010: Data_out <= 16'hA5D7	;
				14'b11100000001011: Data_out <= 16'hA5E0	;
				14'b11100000001100: Data_out <= 16'hA5E9	;
				14'b11100000001101: Data_out <= 16'hA5F2	;
				14'b11100000001110: Data_out <= 16'hA5FB	;
				14'b11100000001111: Data_out <= 16'hA604	;
				14'b11100000010000: Data_out <= 16'hA60D	;
				14'b11100000010001: Data_out <= 16'hA616	;
				14'b11100000010010: Data_out <= 16'hA61F	;
				14'b11100000010011: Data_out <= 16'hA628	;
				14'b11100000010100: Data_out <= 16'hA631	;
				14'b11100000010101: Data_out <= 16'hA63A	;
				14'b11100000010110: Data_out <= 16'hA643	;
				14'b11100000010111: Data_out <= 16'hA64C	;
				14'b11100000011000: Data_out <= 16'hA655	;
				14'b11100000011001: Data_out <= 16'hA65E	;
				14'b11100000011010: Data_out <= 16'hA667	;
				14'b11100000011011: Data_out <= 16'hA66F	;
				14'b11100000011100: Data_out <= 16'hA678	;
				14'b11100000011101: Data_out <= 16'hA681	;
				14'b11100000011110: Data_out <= 16'hA68A	;
				14'b11100000011111: Data_out <= 16'hA693	;
				14'b11100000100000: Data_out <= 16'hA69C	;
				14'b11100000100001: Data_out <= 16'hA6A5	;
				14'b11100000100010: Data_out <= 16'hA6AE	;
				14'b11100000100011: Data_out <= 16'hA6B7	;
				14'b11100000100100: Data_out <= 16'hA6C0	;
				14'b11100000100101: Data_out <= 16'hA6C9	;
				14'b11100000100110: Data_out <= 16'hA6D2	;
				14'b11100000100111: Data_out <= 16'hA6DB	;
				14'b11100000101000: Data_out <= 16'hA6E4	;
				14'b11100000101001: Data_out <= 16'hA6ED	;
				14'b11100000101010: Data_out <= 16'hA6F7	;
				14'b11100000101011: Data_out <= 16'hA700	;
				14'b11100000101100: Data_out <= 16'hA709	;
				14'b11100000101101: Data_out <= 16'hA712	;
				14'b11100000101110: Data_out <= 16'hA71B	;
				14'b11100000101111: Data_out <= 16'hA724	;
				14'b11100000110000: Data_out <= 16'hA72D	;
				14'b11100000110001: Data_out <= 16'hA736	;
				14'b11100000110010: Data_out <= 16'hA73F	;
				14'b11100000110011: Data_out <= 16'hA748	;
				14'b11100000110100: Data_out <= 16'hA751	;
				14'b11100000110101: Data_out <= 16'hA75A	;
				14'b11100000110110: Data_out <= 16'hA763	;
				14'b11100000110111: Data_out <= 16'hA76C	;
				14'b11100000111000: Data_out <= 16'hA775	;
				14'b11100000111001: Data_out <= 16'hA77E	;
				14'b11100000111010: Data_out <= 16'hA787	;
				14'b11100000111011: Data_out <= 16'hA790	;
				14'b11100000111100: Data_out <= 16'hA79A	;
				14'b11100000111101: Data_out <= 16'hA7A3	;
				14'b11100000111110: Data_out <= 16'hA7AC	;
				14'b11100000111111: Data_out <= 16'hA7B5	;
				14'b11100001000000: Data_out <= 16'hA7BE	;
				14'b11100001000001: Data_out <= 16'hA7C7	;
				14'b11100001000010: Data_out <= 16'hA7D0	;
				14'b11100001000011: Data_out <= 16'hA7D9	;
				14'b11100001000100: Data_out <= 16'hA7E2	;
				14'b11100001000101: Data_out <= 16'hA7EB	;
				14'b11100001000110: Data_out <= 16'hA7F5	;
				14'b11100001000111: Data_out <= 16'hA7FE	;
				14'b11100001001000: Data_out <= 16'hA807	;
				14'b11100001001001: Data_out <= 16'hA810	;
				14'b11100001001010: Data_out <= 16'hA819	;
				14'b11100001001011: Data_out <= 16'hA822	;
				14'b11100001001100: Data_out <= 16'hA82B	;
				14'b11100001001101: Data_out <= 16'hA835	;
				14'b11100001001110: Data_out <= 16'hA83E	;
				14'b11100001001111: Data_out <= 16'hA847	;
				14'b11100001010000: Data_out <= 16'hA850	;
				14'b11100001010001: Data_out <= 16'hA859	;
				14'b11100001010010: Data_out <= 16'hA862	;
				14'b11100001010011: Data_out <= 16'hA86B	;
				14'b11100001010100: Data_out <= 16'hA875	;
				14'b11100001010101: Data_out <= 16'hA87E	;
				14'b11100001010110: Data_out <= 16'hA887	;
				14'b11100001010111: Data_out <= 16'hA890	;
				14'b11100001011000: Data_out <= 16'hA899	;
				14'b11100001011001: Data_out <= 16'hA8A2	;
				14'b11100001011010: Data_out <= 16'hA8AC	;
				14'b11100001011011: Data_out <= 16'hA8B5	;
				14'b11100001011100: Data_out <= 16'hA8BE	;
				14'b11100001011101: Data_out <= 16'hA8C7	;
				14'b11100001011110: Data_out <= 16'hA8D0	;
				14'b11100001011111: Data_out <= 16'hA8DA	;
				14'b11100001100000: Data_out <= 16'hA8E3	;
				14'b11100001100001: Data_out <= 16'hA8EC	;
				14'b11100001100010: Data_out <= 16'hA8F5	;
				14'b11100001100011: Data_out <= 16'hA8FE	;
				14'b11100001100100: Data_out <= 16'hA908	;
				14'b11100001100101: Data_out <= 16'hA911	;
				14'b11100001100110: Data_out <= 16'hA91A	;
				14'b11100001100111: Data_out <= 16'hA923	;
				14'b11100001101000: Data_out <= 16'hA92D	;
				14'b11100001101001: Data_out <= 16'hA936	;
				14'b11100001101010: Data_out <= 16'hA93F	;
				14'b11100001101011: Data_out <= 16'hA948	;
				14'b11100001101100: Data_out <= 16'hA952	;
				14'b11100001101101: Data_out <= 16'hA95B	;
				14'b11100001101110: Data_out <= 16'hA964	;
				14'b11100001101111: Data_out <= 16'hA96D	;
				14'b11100001110000: Data_out <= 16'hA977	;
				14'b11100001110001: Data_out <= 16'hA980	;
				14'b11100001110010: Data_out <= 16'hA989	;
				14'b11100001110011: Data_out <= 16'hA992	;
				14'b11100001110100: Data_out <= 16'hA99C	;
				14'b11100001110101: Data_out <= 16'hA9A5	;
				14'b11100001110110: Data_out <= 16'hA9AE	;
				14'b11100001110111: Data_out <= 16'hA9B7	;
				14'b11100001111000: Data_out <= 16'hA9C1	;
				14'b11100001111001: Data_out <= 16'hA9CA	;
				14'b11100001111010: Data_out <= 16'hA9D3	;
				14'b11100001111011: Data_out <= 16'hA9DD	;
				14'b11100001111100: Data_out <= 16'hA9E6	;
				14'b11100001111101: Data_out <= 16'hA9EF	;
				14'b11100001111110: Data_out <= 16'hA9F9	;
				14'b11100001111111: Data_out <= 16'hAA02	;
				14'b11100010000000: Data_out <= 16'hAA0B	;
				14'b11100010000001: Data_out <= 16'hAA14	;
				14'b11100010000010: Data_out <= 16'hAA1E	;
				14'b11100010000011: Data_out <= 16'hAA27	;
				14'b11100010000100: Data_out <= 16'hAA30	;
				14'b11100010000101: Data_out <= 16'hAA3A	;
				14'b11100010000110: Data_out <= 16'hAA43	;
				14'b11100010000111: Data_out <= 16'hAA4C	;
				14'b11100010001000: Data_out <= 16'hAA56	;
				14'b11100010001001: Data_out <= 16'hAA5F	;
				14'b11100010001010: Data_out <= 16'hAA68	;
				14'b11100010001011: Data_out <= 16'hAA72	;
				14'b11100010001100: Data_out <= 16'hAA7B	;
				14'b11100010001101: Data_out <= 16'hAA84	;
				14'b11100010001110: Data_out <= 16'hAA8E	;
				14'b11100010001111: Data_out <= 16'hAA97	;
				14'b11100010010000: Data_out <= 16'hAAA1	;
				14'b11100010010001: Data_out <= 16'hAAAA	;
				14'b11100010010010: Data_out <= 16'hAAB3	;
				14'b11100010010011: Data_out <= 16'hAABD	;
				14'b11100010010100: Data_out <= 16'hAAC6	;
				14'b11100010010101: Data_out <= 16'hAACF	;
				14'b11100010010110: Data_out <= 16'hAAD9	;
				14'b11100010010111: Data_out <= 16'hAAE2	;
				14'b11100010011000: Data_out <= 16'hAAEC	;
				14'b11100010011001: Data_out <= 16'hAAF5	;
				14'b11100010011010: Data_out <= 16'hAAFE	;
				14'b11100010011011: Data_out <= 16'hAB08	;
				14'b11100010011100: Data_out <= 16'hAB11	;
				14'b11100010011101: Data_out <= 16'hAB1A	;
				14'b11100010011110: Data_out <= 16'hAB24	;
				14'b11100010011111: Data_out <= 16'hAB2D	;
				14'b11100010100000: Data_out <= 16'hAB37	;
				14'b11100010100001: Data_out <= 16'hAB40	;
				14'b11100010100010: Data_out <= 16'hAB4A	;
				14'b11100010100011: Data_out <= 16'hAB53	;
				14'b11100010100100: Data_out <= 16'hAB5C	;
				14'b11100010100101: Data_out <= 16'hAB66	;
				14'b11100010100110: Data_out <= 16'hAB6F	;
				14'b11100010100111: Data_out <= 16'hAB79	;
				14'b11100010101000: Data_out <= 16'hAB82	;
				14'b11100010101001: Data_out <= 16'hAB8C	;
				14'b11100010101010: Data_out <= 16'hAB95	;
				14'b11100010101011: Data_out <= 16'hAB9E	;
				14'b11100010101100: Data_out <= 16'hABA8	;
				14'b11100010101101: Data_out <= 16'hABB1	;
				14'b11100010101110: Data_out <= 16'hABBB	;
				14'b11100010101111: Data_out <= 16'hABC4	;
				14'b11100010110000: Data_out <= 16'hABCE	;
				14'b11100010110001: Data_out <= 16'hABD7	;
				14'b11100010110010: Data_out <= 16'hABE1	;
				14'b11100010110011: Data_out <= 16'hABEA	;
				14'b11100010110100: Data_out <= 16'hABF4	;
				14'b11100010110101: Data_out <= 16'hABFD	;
				14'b11100010110110: Data_out <= 16'hAC07	;
				14'b11100010110111: Data_out <= 16'hAC10	;
				14'b11100010111000: Data_out <= 16'hAC1A	;
				14'b11100010111001: Data_out <= 16'hAC23	;
				14'b11100010111010: Data_out <= 16'hAC2D	;
				14'b11100010111011: Data_out <= 16'hAC36	;
				14'b11100010111100: Data_out <= 16'hAC40	;
				14'b11100010111101: Data_out <= 16'hAC49	;
				14'b11100010111110: Data_out <= 16'hAC53	;
				14'b11100010111111: Data_out <= 16'hAC5C	;
				14'b11100011000000: Data_out <= 16'hAC66	;
				14'b11100011000001: Data_out <= 16'hAC6F	;
				14'b11100011000010: Data_out <= 16'hAC79	;
				14'b11100011000011: Data_out <= 16'hAC82	;
				14'b11100011000100: Data_out <= 16'hAC8C	;
				14'b11100011000101: Data_out <= 16'hAC95	;
				14'b11100011000110: Data_out <= 16'hAC9F	;
				14'b11100011000111: Data_out <= 16'hACA8	;
				14'b11100011001000: Data_out <= 16'hACB2	;
				14'b11100011001001: Data_out <= 16'hACBB	;
				14'b11100011001010: Data_out <= 16'hACC5	;
				14'b11100011001011: Data_out <= 16'hACCE	;
				14'b11100011001100: Data_out <= 16'hACD8	;
				14'b11100011001101: Data_out <= 16'hACE2	;
				14'b11100011001110: Data_out <= 16'hACEB	;
				14'b11100011001111: Data_out <= 16'hACF5	;
				14'b11100011010000: Data_out <= 16'hACFE	;
				14'b11100011010001: Data_out <= 16'hAD08	;
				14'b11100011010010: Data_out <= 16'hAD11	;
				14'b11100011010011: Data_out <= 16'hAD1B	;
				14'b11100011010100: Data_out <= 16'hAD25	;
				14'b11100011010101: Data_out <= 16'hAD2E	;
				14'b11100011010110: Data_out <= 16'hAD38	;
				14'b11100011010111: Data_out <= 16'hAD41	;
				14'b11100011011000: Data_out <= 16'hAD4B	;
				14'b11100011011001: Data_out <= 16'hAD54	;
				14'b11100011011010: Data_out <= 16'hAD5E	;
				14'b11100011011011: Data_out <= 16'hAD68	;
				14'b11100011011100: Data_out <= 16'hAD71	;
				14'b11100011011101: Data_out <= 16'hAD7B	;
				14'b11100011011110: Data_out <= 16'hAD84	;
				14'b11100011011111: Data_out <= 16'hAD8E	;
				14'b11100011100000: Data_out <= 16'hAD98	;
				14'b11100011100001: Data_out <= 16'hADA1	;
				14'b11100011100010: Data_out <= 16'hADAB	;
				14'b11100011100011: Data_out <= 16'hADB5	;
				14'b11100011100100: Data_out <= 16'hADBE	;
				14'b11100011100101: Data_out <= 16'hADC8	;
				14'b11100011100110: Data_out <= 16'hADD1	;
				14'b11100011100111: Data_out <= 16'hADDB	;
				14'b11100011101000: Data_out <= 16'hADE5	;
				14'b11100011101001: Data_out <= 16'hADEE	;
				14'b11100011101010: Data_out <= 16'hADF8	;
				14'b11100011101011: Data_out <= 16'hAE02	;
				14'b11100011101100: Data_out <= 16'hAE0B	;
				14'b11100011101101: Data_out <= 16'hAE15	;
				14'b11100011101110: Data_out <= 16'hAE1F	;
				14'b11100011101111: Data_out <= 16'hAE28	;
				14'b11100011110000: Data_out <= 16'hAE32	;
				14'b11100011110001: Data_out <= 16'hAE3C	;
				14'b11100011110010: Data_out <= 16'hAE45	;
				14'b11100011110011: Data_out <= 16'hAE4F	;
				14'b11100011110100: Data_out <= 16'hAE59	;
				14'b11100011110101: Data_out <= 16'hAE62	;
				14'b11100011110110: Data_out <= 16'hAE6C	;
				14'b11100011110111: Data_out <= 16'hAE76	;
				14'b11100011111000: Data_out <= 16'hAE7F	;
				14'b11100011111001: Data_out <= 16'hAE89	;
				14'b11100011111010: Data_out <= 16'hAE93	;
				14'b11100011111011: Data_out <= 16'hAE9C	;
				14'b11100011111100: Data_out <= 16'hAEA6	;
				14'b11100011111101: Data_out <= 16'hAEB0	;
				14'b11100011111110: Data_out <= 16'hAEBA	;
				14'b11100011111111: Data_out <= 16'hAEC3	;
				14'b11100100000000: Data_out <= 16'hAECD	;
				14'b11100100000001: Data_out <= 16'hAED7	;
				14'b11100100000010: Data_out <= 16'hAEE0	;
				14'b11100100000011: Data_out <= 16'hAEEA	;
				14'b11100100000100: Data_out <= 16'hAEF4	;
				14'b11100100000101: Data_out <= 16'hAEFE	;
				14'b11100100000110: Data_out <= 16'hAF07	;
				14'b11100100000111: Data_out <= 16'hAF11	;
				14'b11100100001000: Data_out <= 16'hAF1B	;
				14'b11100100001001: Data_out <= 16'hAF24	;
				14'b11100100001010: Data_out <= 16'hAF2E	;
				14'b11100100001011: Data_out <= 16'hAF38	;
				14'b11100100001100: Data_out <= 16'hAF42	;
				14'b11100100001101: Data_out <= 16'hAF4B	;
				14'b11100100001110: Data_out <= 16'hAF55	;
				14'b11100100001111: Data_out <= 16'hAF5F	;
				14'b11100100010000: Data_out <= 16'hAF69	;
				14'b11100100010001: Data_out <= 16'hAF73	;
				14'b11100100010010: Data_out <= 16'hAF7C	;
				14'b11100100010011: Data_out <= 16'hAF86	;
				14'b11100100010100: Data_out <= 16'hAF90	;
				14'b11100100010101: Data_out <= 16'hAF9A	;
				14'b11100100010110: Data_out <= 16'hAFA3	;
				14'b11100100010111: Data_out <= 16'hAFAD	;
				14'b11100100011000: Data_out <= 16'hAFB7	;
				14'b11100100011001: Data_out <= 16'hAFC1	;
				14'b11100100011010: Data_out <= 16'hAFCB	;
				14'b11100100011011: Data_out <= 16'hAFD4	;
				14'b11100100011100: Data_out <= 16'hAFDE	;
				14'b11100100011101: Data_out <= 16'hAFE8	;
				14'b11100100011110: Data_out <= 16'hAFF2	;
				14'b11100100011111: Data_out <= 16'hAFFC	;
				14'b11100100100000: Data_out <= 16'hB005	;
				14'b11100100100001: Data_out <= 16'hB00F	;
				14'b11100100100010: Data_out <= 16'hB019	;
				14'b11100100100011: Data_out <= 16'hB023	;
				14'b11100100100100: Data_out <= 16'hB02D	;
				14'b11100100100101: Data_out <= 16'hB036	;
				14'b11100100100110: Data_out <= 16'hB040	;
				14'b11100100100111: Data_out <= 16'hB04A	;
				14'b11100100101000: Data_out <= 16'hB054	;
				14'b11100100101001: Data_out <= 16'hB05E	;
				14'b11100100101010: Data_out <= 16'hB068	;
				14'b11100100101011: Data_out <= 16'hB071	;
				14'b11100100101100: Data_out <= 16'hB07B	;
				14'b11100100101101: Data_out <= 16'hB085	;
				14'b11100100101110: Data_out <= 16'hB08F	;
				14'b11100100101111: Data_out <= 16'hB099	;
				14'b11100100110000: Data_out <= 16'hB0A3	;
				14'b11100100110001: Data_out <= 16'hB0AD	;
				14'b11100100110010: Data_out <= 16'hB0B6	;
				14'b11100100110011: Data_out <= 16'hB0C0	;
				14'b11100100110100: Data_out <= 16'hB0CA	;
				14'b11100100110101: Data_out <= 16'hB0D4	;
				14'b11100100110110: Data_out <= 16'hB0DE	;
				14'b11100100110111: Data_out <= 16'hB0E8	;
				14'b11100100111000: Data_out <= 16'hB0F2	;
				14'b11100100111001: Data_out <= 16'hB0FC	;
				14'b11100100111010: Data_out <= 16'hB105	;
				14'b11100100111011: Data_out <= 16'hB10F	;
				14'b11100100111100: Data_out <= 16'hB119	;
				14'b11100100111101: Data_out <= 16'hB123	;
				14'b11100100111110: Data_out <= 16'hB12D	;
				14'b11100100111111: Data_out <= 16'hB137	;
				14'b11100101000000: Data_out <= 16'hB141	;
				14'b11100101000001: Data_out <= 16'hB14B	;
				14'b11100101000010: Data_out <= 16'hB155	;
				14'b11100101000011: Data_out <= 16'hB15F	;
				14'b11100101000100: Data_out <= 16'hB168	;
				14'b11100101000101: Data_out <= 16'hB172	;
				14'b11100101000110: Data_out <= 16'hB17C	;
				14'b11100101000111: Data_out <= 16'hB186	;
				14'b11100101001000: Data_out <= 16'hB190	;
				14'b11100101001001: Data_out <= 16'hB19A	;
				14'b11100101001010: Data_out <= 16'hB1A4	;
				14'b11100101001011: Data_out <= 16'hB1AE	;
				14'b11100101001100: Data_out <= 16'hB1B8	;
				14'b11100101001101: Data_out <= 16'hB1C2	;
				14'b11100101001110: Data_out <= 16'hB1CC	;
				14'b11100101001111: Data_out <= 16'hB1D6	;
				14'b11100101010000: Data_out <= 16'hB1E0	;
				14'b11100101010001: Data_out <= 16'hB1EA	;
				14'b11100101010010: Data_out <= 16'hB1F4	;
				14'b11100101010011: Data_out <= 16'hB1FE	;
				14'b11100101010100: Data_out <= 16'hB208	;
				14'b11100101010101: Data_out <= 16'hB211	;
				14'b11100101010110: Data_out <= 16'hB21B	;
				14'b11100101010111: Data_out <= 16'hB225	;
				14'b11100101011000: Data_out <= 16'hB22F	;
				14'b11100101011001: Data_out <= 16'hB239	;
				14'b11100101011010: Data_out <= 16'hB243	;
				14'b11100101011011: Data_out <= 16'hB24D	;
				14'b11100101011100: Data_out <= 16'hB257	;
				14'b11100101011101: Data_out <= 16'hB261	;
				14'b11100101011110: Data_out <= 16'hB26B	;
				14'b11100101011111: Data_out <= 16'hB275	;
				14'b11100101100000: Data_out <= 16'hB27F	;
				14'b11100101100001: Data_out <= 16'hB289	;
				14'b11100101100010: Data_out <= 16'hB293	;
				14'b11100101100011: Data_out <= 16'hB29D	;
				14'b11100101100100: Data_out <= 16'hB2A7	;
				14'b11100101100101: Data_out <= 16'hB2B1	;
				14'b11100101100110: Data_out <= 16'hB2BB	;
				14'b11100101100111: Data_out <= 16'hB2C5	;
				14'b11100101101000: Data_out <= 16'hB2CF	;
				14'b11100101101001: Data_out <= 16'hB2D9	;
				14'b11100101101010: Data_out <= 16'hB2E3	;
				14'b11100101101011: Data_out <= 16'hB2EE	;
				14'b11100101101100: Data_out <= 16'hB2F8	;
				14'b11100101101101: Data_out <= 16'hB302	;
				14'b11100101101110: Data_out <= 16'hB30C	;
				14'b11100101101111: Data_out <= 16'hB316	;
				14'b11100101110000: Data_out <= 16'hB320	;
				14'b11100101110001: Data_out <= 16'hB32A	;
				14'b11100101110010: Data_out <= 16'hB334	;
				14'b11100101110011: Data_out <= 16'hB33E	;
				14'b11100101110100: Data_out <= 16'hB348	;
				14'b11100101110101: Data_out <= 16'hB352	;
				14'b11100101110110: Data_out <= 16'hB35C	;
				14'b11100101110111: Data_out <= 16'hB366	;
				14'b11100101111000: Data_out <= 16'hB370	;
				14'b11100101111001: Data_out <= 16'hB37A	;
				14'b11100101111010: Data_out <= 16'hB384	;
				14'b11100101111011: Data_out <= 16'hB38E	;
				14'b11100101111100: Data_out <= 16'hB398	;
				14'b11100101111101: Data_out <= 16'hB3A3	;
				14'b11100101111110: Data_out <= 16'hB3AD	;
				14'b11100101111111: Data_out <= 16'hB3B7	;
				14'b11100110000000: Data_out <= 16'hB3C1	;
				14'b11100110000001: Data_out <= 16'hB3CB	;
				14'b11100110000010: Data_out <= 16'hB3D5	;
				14'b11100110000011: Data_out <= 16'hB3DF	;
				14'b11100110000100: Data_out <= 16'hB3E9	;
				14'b11100110000101: Data_out <= 16'hB3F3	;
				14'b11100110000110: Data_out <= 16'hB3FD	;
				14'b11100110000111: Data_out <= 16'hB408	;
				14'b11100110001000: Data_out <= 16'hB412	;
				14'b11100110001001: Data_out <= 16'hB41C	;
				14'b11100110001010: Data_out <= 16'hB426	;
				14'b11100110001011: Data_out <= 16'hB430	;
				14'b11100110001100: Data_out <= 16'hB43A	;
				14'b11100110001101: Data_out <= 16'hB444	;
				14'b11100110001110: Data_out <= 16'hB44E	;
				14'b11100110001111: Data_out <= 16'hB459	;
				14'b11100110010000: Data_out <= 16'hB463	;
				14'b11100110010001: Data_out <= 16'hB46D	;
				14'b11100110010010: Data_out <= 16'hB477	;
				14'b11100110010011: Data_out <= 16'hB481	;
				14'b11100110010100: Data_out <= 16'hB48B	;
				14'b11100110010101: Data_out <= 16'hB495	;
				14'b11100110010110: Data_out <= 16'hB4A0	;
				14'b11100110010111: Data_out <= 16'hB4AA	;
				14'b11100110011000: Data_out <= 16'hB4B4	;
				14'b11100110011001: Data_out <= 16'hB4BE	;
				14'b11100110011010: Data_out <= 16'hB4C8	;
				14'b11100110011011: Data_out <= 16'hB4D2	;
				14'b11100110011100: Data_out <= 16'hB4DD	;
				14'b11100110011101: Data_out <= 16'hB4E7	;
				14'b11100110011110: Data_out <= 16'hB4F1	;
				14'b11100110011111: Data_out <= 16'hB4FB	;
				14'b11100110100000: Data_out <= 16'hB505	;
				14'b11100110100001: Data_out <= 16'hB50F	;
				14'b11100110100010: Data_out <= 16'hB51A	;
				14'b11100110100011: Data_out <= 16'hB524	;
				14'b11100110100100: Data_out <= 16'hB52E	;
				14'b11100110100101: Data_out <= 16'hB538	;
				14'b11100110100110: Data_out <= 16'hB542	;
				14'b11100110100111: Data_out <= 16'hB54D	;
				14'b11100110101000: Data_out <= 16'hB557	;
				14'b11100110101001: Data_out <= 16'hB561	;
				14'b11100110101010: Data_out <= 16'hB56B	;
				14'b11100110101011: Data_out <= 16'hB575	;
				14'b11100110101100: Data_out <= 16'hB580	;
				14'b11100110101101: Data_out <= 16'hB58A	;
				14'b11100110101110: Data_out <= 16'hB594	;
				14'b11100110101111: Data_out <= 16'hB59E	;
				14'b11100110110000: Data_out <= 16'hB5A9	;
				14'b11100110110001: Data_out <= 16'hB5B3	;
				14'b11100110110010: Data_out <= 16'hB5BD	;
				14'b11100110110011: Data_out <= 16'hB5C7	;
				14'b11100110110100: Data_out <= 16'hB5D2	;
				14'b11100110110101: Data_out <= 16'hB5DC	;
				14'b11100110110110: Data_out <= 16'hB5E6	;
				14'b11100110110111: Data_out <= 16'hB5F0	;
				14'b11100110111000: Data_out <= 16'hB5FA	;
				14'b11100110111001: Data_out <= 16'hB605	;
				14'b11100110111010: Data_out <= 16'hB60F	;
				14'b11100110111011: Data_out <= 16'hB619	;
				14'b11100110111100: Data_out <= 16'hB624	;
				14'b11100110111101: Data_out <= 16'hB62E	;
				14'b11100110111110: Data_out <= 16'hB638	;
				14'b11100110111111: Data_out <= 16'hB642	;
				14'b11100111000000: Data_out <= 16'hB64D	;
				14'b11100111000001: Data_out <= 16'hB657	;
				14'b11100111000010: Data_out <= 16'hB661	;
				14'b11100111000011: Data_out <= 16'hB66B	;
				14'b11100111000100: Data_out <= 16'hB676	;
				14'b11100111000101: Data_out <= 16'hB680	;
				14'b11100111000110: Data_out <= 16'hB68A	;
				14'b11100111000111: Data_out <= 16'hB695	;
				14'b11100111001000: Data_out <= 16'hB69F	;
				14'b11100111001001: Data_out <= 16'hB6A9	;
				14'b11100111001010: Data_out <= 16'hB6B3	;
				14'b11100111001011: Data_out <= 16'hB6BE	;
				14'b11100111001100: Data_out <= 16'hB6C8	;
				14'b11100111001101: Data_out <= 16'hB6D2	;
				14'b11100111001110: Data_out <= 16'hB6DD	;
				14'b11100111001111: Data_out <= 16'hB6E7	;
				14'b11100111010000: Data_out <= 16'hB6F1	;
				14'b11100111010001: Data_out <= 16'hB6FC	;
				14'b11100111010010: Data_out <= 16'hB706	;
				14'b11100111010011: Data_out <= 16'hB710	;
				14'b11100111010100: Data_out <= 16'hB71B	;
				14'b11100111010101: Data_out <= 16'hB725	;
				14'b11100111010110: Data_out <= 16'hB72F	;
				14'b11100111010111: Data_out <= 16'hB73A	;
				14'b11100111011000: Data_out <= 16'hB744	;
				14'b11100111011001: Data_out <= 16'hB74E	;
				14'b11100111011010: Data_out <= 16'hB759	;
				14'b11100111011011: Data_out <= 16'hB763	;
				14'b11100111011100: Data_out <= 16'hB76D	;
				14'b11100111011101: Data_out <= 16'hB778	;
				14'b11100111011110: Data_out <= 16'hB782	;
				14'b11100111011111: Data_out <= 16'hB78C	;
				14'b11100111100000: Data_out <= 16'hB797	;
				14'b11100111100001: Data_out <= 16'hB7A1	;
				14'b11100111100010: Data_out <= 16'hB7AB	;
				14'b11100111100011: Data_out <= 16'hB7B6	;
				14'b11100111100100: Data_out <= 16'hB7C0	;
				14'b11100111100101: Data_out <= 16'hB7CB	;
				14'b11100111100110: Data_out <= 16'hB7D5	;
				14'b11100111100111: Data_out <= 16'hB7DF	;
				14'b11100111101000: Data_out <= 16'hB7EA	;
				14'b11100111101001: Data_out <= 16'hB7F4	;
				14'b11100111101010: Data_out <= 16'hB7FF	;
				14'b11100111101011: Data_out <= 16'hB809	;
				14'b11100111101100: Data_out <= 16'hB813	;
				14'b11100111101101: Data_out <= 16'hB81E	;
				14'b11100111101110: Data_out <= 16'hB828	;
				14'b11100111101111: Data_out <= 16'hB832	;
				14'b11100111110000: Data_out <= 16'hB83D	;
				14'b11100111110001: Data_out <= 16'hB847	;
				14'b11100111110010: Data_out <= 16'hB852	;
				14'b11100111110011: Data_out <= 16'hB85C	;
				14'b11100111110100: Data_out <= 16'hB867	;
				14'b11100111110101: Data_out <= 16'hB871	;
				14'b11100111110110: Data_out <= 16'hB87B	;
				14'b11100111110111: Data_out <= 16'hB886	;
				14'b11100111111000: Data_out <= 16'hB890	;
				14'b11100111111001: Data_out <= 16'hB89B	;
				14'b11100111111010: Data_out <= 16'hB8A5	;
				14'b11100111111011: Data_out <= 16'hB8B0	;
				14'b11100111111100: Data_out <= 16'hB8BA	;
				14'b11100111111101: Data_out <= 16'hB8C4	;
				14'b11100111111110: Data_out <= 16'hB8CF	;
				14'b11100111111111: Data_out <= 16'hB8D9	;
				14'b11101000000000: Data_out <= 16'hB8E4	;
				14'b11101000000001: Data_out <= 16'hB8EE	;
				14'b11101000000010: Data_out <= 16'hB8F9	;
				14'b11101000000011: Data_out <= 16'hB903	;
				14'b11101000000100: Data_out <= 16'hB90E	;
				14'b11101000000101: Data_out <= 16'hB918	;
				14'b11101000000110: Data_out <= 16'hB922	;
				14'b11101000000111: Data_out <= 16'hB92D	;
				14'b11101000001000: Data_out <= 16'hB937	;
				14'b11101000001001: Data_out <= 16'hB942	;
				14'b11101000001010: Data_out <= 16'hB94C	;
				14'b11101000001011: Data_out <= 16'hB957	;
				14'b11101000001100: Data_out <= 16'hB961	;
				14'b11101000001101: Data_out <= 16'hB96C	;
				14'b11101000001110: Data_out <= 16'hB976	;
				14'b11101000001111: Data_out <= 16'hB981	;
				14'b11101000010000: Data_out <= 16'hB98B	;
				14'b11101000010001: Data_out <= 16'hB996	;
				14'b11101000010010: Data_out <= 16'hB9A0	;
				14'b11101000010011: Data_out <= 16'hB9AB	;
				14'b11101000010100: Data_out <= 16'hB9B5	;
				14'b11101000010101: Data_out <= 16'hB9C0	;
				14'b11101000010110: Data_out <= 16'hB9CA	;
				14'b11101000010111: Data_out <= 16'hB9D5	;
				14'b11101000011000: Data_out <= 16'hB9DF	;
				14'b11101000011001: Data_out <= 16'hB9EA	;
				14'b11101000011010: Data_out <= 16'hB9F4	;
				14'b11101000011011: Data_out <= 16'hB9FF	;
				14'b11101000011100: Data_out <= 16'hBA09	;
				14'b11101000011101: Data_out <= 16'hBA14	;
				14'b11101000011110: Data_out <= 16'hBA1E	;
				14'b11101000011111: Data_out <= 16'hBA29	;
				14'b11101000100000: Data_out <= 16'hBA33	;
				14'b11101000100001: Data_out <= 16'hBA3E	;
				14'b11101000100010: Data_out <= 16'hBA49	;
				14'b11101000100011: Data_out <= 16'hBA53	;
				14'b11101000100100: Data_out <= 16'hBA5E	;
				14'b11101000100101: Data_out <= 16'hBA68	;
				14'b11101000100110: Data_out <= 16'hBA73	;
				14'b11101000100111: Data_out <= 16'hBA7D	;
				14'b11101000101000: Data_out <= 16'hBA88	;
				14'b11101000101001: Data_out <= 16'hBA92	;
				14'b11101000101010: Data_out <= 16'hBA9D	;
				14'b11101000101011: Data_out <= 16'hBAA7	;
				14'b11101000101100: Data_out <= 16'hBAB2	;
				14'b11101000101101: Data_out <= 16'hBABD	;
				14'b11101000101110: Data_out <= 16'hBAC7	;
				14'b11101000101111: Data_out <= 16'hBAD2	;
				14'b11101000110000: Data_out <= 16'hBADC	;
				14'b11101000110001: Data_out <= 16'hBAE7	;
				14'b11101000110010: Data_out <= 16'hBAF1	;
				14'b11101000110011: Data_out <= 16'hBAFC	;
				14'b11101000110100: Data_out <= 16'hBB07	;
				14'b11101000110101: Data_out <= 16'hBB11	;
				14'b11101000110110: Data_out <= 16'hBB1C	;
				14'b11101000110111: Data_out <= 16'hBB26	;
				14'b11101000111000: Data_out <= 16'hBB31	;
				14'b11101000111001: Data_out <= 16'hBB3C	;
				14'b11101000111010: Data_out <= 16'hBB46	;
				14'b11101000111011: Data_out <= 16'hBB51	;
				14'b11101000111100: Data_out <= 16'hBB5B	;
				14'b11101000111101: Data_out <= 16'hBB66	;
				14'b11101000111110: Data_out <= 16'hBB71	;
				14'b11101000111111: Data_out <= 16'hBB7B	;
				14'b11101001000000: Data_out <= 16'hBB86	;
				14'b11101001000001: Data_out <= 16'hBB90	;
				14'b11101001000010: Data_out <= 16'hBB9B	;
				14'b11101001000011: Data_out <= 16'hBBA6	;
				14'b11101001000100: Data_out <= 16'hBBB0	;
				14'b11101001000101: Data_out <= 16'hBBBB	;
				14'b11101001000110: Data_out <= 16'hBBC6	;
				14'b11101001000111: Data_out <= 16'hBBD0	;
				14'b11101001001000: Data_out <= 16'hBBDB	;
				14'b11101001001001: Data_out <= 16'hBBE5	;
				14'b11101001001010: Data_out <= 16'hBBF0	;
				14'b11101001001011: Data_out <= 16'hBBFB	;
				14'b11101001001100: Data_out <= 16'hBC05	;
				14'b11101001001101: Data_out <= 16'hBC10	;
				14'b11101001001110: Data_out <= 16'hBC1B	;
				14'b11101001001111: Data_out <= 16'hBC25	;
				14'b11101001010000: Data_out <= 16'hBC30	;
				14'b11101001010001: Data_out <= 16'hBC3B	;
				14'b11101001010010: Data_out <= 16'hBC45	;
				14'b11101001010011: Data_out <= 16'hBC50	;
				14'b11101001010100: Data_out <= 16'hBC5B	;
				14'b11101001010101: Data_out <= 16'hBC65	;
				14'b11101001010110: Data_out <= 16'hBC70	;
				14'b11101001010111: Data_out <= 16'hBC7B	;
				14'b11101001011000: Data_out <= 16'hBC85	;
				14'b11101001011001: Data_out <= 16'hBC90	;
				14'b11101001011010: Data_out <= 16'hBC9B	;
				14'b11101001011011: Data_out <= 16'hBCA5	;
				14'b11101001011100: Data_out <= 16'hBCB0	;
				14'b11101001011101: Data_out <= 16'hBCBB	;
				14'b11101001011110: Data_out <= 16'hBCC5	;
				14'b11101001011111: Data_out <= 16'hBCD0	;
				14'b11101001100000: Data_out <= 16'hBCDB	;
				14'b11101001100001: Data_out <= 16'hBCE6	;
				14'b11101001100010: Data_out <= 16'hBCF0	;
				14'b11101001100011: Data_out <= 16'hBCFB	;
				14'b11101001100100: Data_out <= 16'hBD06	;
				14'b11101001100101: Data_out <= 16'hBD10	;
				14'b11101001100110: Data_out <= 16'hBD1B	;
				14'b11101001100111: Data_out <= 16'hBD26	;
				14'b11101001101000: Data_out <= 16'hBD31	;
				14'b11101001101001: Data_out <= 16'hBD3B	;
				14'b11101001101010: Data_out <= 16'hBD46	;
				14'b11101001101011: Data_out <= 16'hBD51	;
				14'b11101001101100: Data_out <= 16'hBD5B	;
				14'b11101001101101: Data_out <= 16'hBD66	;
				14'b11101001101110: Data_out <= 16'hBD71	;
				14'b11101001101111: Data_out <= 16'hBD7C	;
				14'b11101001110000: Data_out <= 16'hBD86	;
				14'b11101001110001: Data_out <= 16'hBD91	;
				14'b11101001110010: Data_out <= 16'hBD9C	;
				14'b11101001110011: Data_out <= 16'hBDA7	;
				14'b11101001110100: Data_out <= 16'hBDB1	;
				14'b11101001110101: Data_out <= 16'hBDBC	;
				14'b11101001110110: Data_out <= 16'hBDC7	;
				14'b11101001110111: Data_out <= 16'hBDD2	;
				14'b11101001111000: Data_out <= 16'hBDDC	;
				14'b11101001111001: Data_out <= 16'hBDE7	;
				14'b11101001111010: Data_out <= 16'hBDF2	;
				14'b11101001111011: Data_out <= 16'hBDFD	;
				14'b11101001111100: Data_out <= 16'hBE07	;
				14'b11101001111101: Data_out <= 16'hBE12	;
				14'b11101001111110: Data_out <= 16'hBE1D	;
				14'b11101001111111: Data_out <= 16'hBE28	;
				14'b11101010000000: Data_out <= 16'hBE32	;
				14'b11101010000001: Data_out <= 16'hBE3D	;
				14'b11101010000010: Data_out <= 16'hBE48	;
				14'b11101010000011: Data_out <= 16'hBE53	;
				14'b11101010000100: Data_out <= 16'hBE5E	;
				14'b11101010000101: Data_out <= 16'hBE68	;
				14'b11101010000110: Data_out <= 16'hBE73	;
				14'b11101010000111: Data_out <= 16'hBE7E	;
				14'b11101010001000: Data_out <= 16'hBE89	;
				14'b11101010001001: Data_out <= 16'hBE94	;
				14'b11101010001010: Data_out <= 16'hBE9E	;
				14'b11101010001011: Data_out <= 16'hBEA9	;
				14'b11101010001100: Data_out <= 16'hBEB4	;
				14'b11101010001101: Data_out <= 16'hBEBF	;
				14'b11101010001110: Data_out <= 16'hBECA	;
				14'b11101010001111: Data_out <= 16'hBED4	;
				14'b11101010010000: Data_out <= 16'hBEDF	;
				14'b11101010010001: Data_out <= 16'hBEEA	;
				14'b11101010010010: Data_out <= 16'hBEF5	;
				14'b11101010010011: Data_out <= 16'hBF00	;
				14'b11101010010100: Data_out <= 16'hBF0B	;
				14'b11101010010101: Data_out <= 16'hBF15	;
				14'b11101010010110: Data_out <= 16'hBF20	;
				14'b11101010010111: Data_out <= 16'hBF2B	;
				14'b11101010011000: Data_out <= 16'hBF36	;
				14'b11101010011001: Data_out <= 16'hBF41	;
				14'b11101010011010: Data_out <= 16'hBF4C	;
				14'b11101010011011: Data_out <= 16'hBF56	;
				14'b11101010011100: Data_out <= 16'hBF61	;
				14'b11101010011101: Data_out <= 16'hBF6C	;
				14'b11101010011110: Data_out <= 16'hBF77	;
				14'b11101010011111: Data_out <= 16'hBF82	;
				14'b11101010100000: Data_out <= 16'hBF8D	;
				14'b11101010100001: Data_out <= 16'hBF98	;
				14'b11101010100010: Data_out <= 16'hBFA2	;
				14'b11101010100011: Data_out <= 16'hBFAD	;
				14'b11101010100100: Data_out <= 16'hBFB8	;
				14'b11101010100101: Data_out <= 16'hBFC3	;
				14'b11101010100110: Data_out <= 16'hBFCE	;
				14'b11101010100111: Data_out <= 16'hBFD9	;
				14'b11101010101000: Data_out <= 16'hBFE4	;
				14'b11101010101001: Data_out <= 16'hBFEE	;
				14'b11101010101010: Data_out <= 16'hBFF9	;
				14'b11101010101011: Data_out <= 16'hC004	;
				14'b11101010101100: Data_out <= 16'hC00F	;
				14'b11101010101101: Data_out <= 16'hC01A	;
				14'b11101010101110: Data_out <= 16'hC025	;
				14'b11101010101111: Data_out <= 16'hC030	;
				14'b11101010110000: Data_out <= 16'hC03B	;
				14'b11101010110001: Data_out <= 16'hC046	;
				14'b11101010110010: Data_out <= 16'hC050	;
				14'b11101010110011: Data_out <= 16'hC05B	;
				14'b11101010110100: Data_out <= 16'hC066	;
				14'b11101010110101: Data_out <= 16'hC071	;
				14'b11101010110110: Data_out <= 16'hC07C	;
				14'b11101010110111: Data_out <= 16'hC087	;
				14'b11101010111000: Data_out <= 16'hC092	;
				14'b11101010111001: Data_out <= 16'hC09D	;
				14'b11101010111010: Data_out <= 16'hC0A8	;
				14'b11101010111011: Data_out <= 16'hC0B3	;
				14'b11101010111100: Data_out <= 16'hC0BE	;
				14'b11101010111101: Data_out <= 16'hC0C9	;
				14'b11101010111110: Data_out <= 16'hC0D3	;
				14'b11101010111111: Data_out <= 16'hC0DE	;
				14'b11101011000000: Data_out <= 16'hC0E9	;
				14'b11101011000001: Data_out <= 16'hC0F4	;
				14'b11101011000010: Data_out <= 16'hC0FF	;
				14'b11101011000011: Data_out <= 16'hC10A	;
				14'b11101011000100: Data_out <= 16'hC115	;
				14'b11101011000101: Data_out <= 16'hC120	;
				14'b11101011000110: Data_out <= 16'hC12B	;
				14'b11101011000111: Data_out <= 16'hC136	;
				14'b11101011001000: Data_out <= 16'hC141	;
				14'b11101011001001: Data_out <= 16'hC14C	;
				14'b11101011001010: Data_out <= 16'hC157	;
				14'b11101011001011: Data_out <= 16'hC162	;
				14'b11101011001100: Data_out <= 16'hC16D	;
				14'b11101011001101: Data_out <= 16'hC178	;
				14'b11101011001110: Data_out <= 16'hC183	;
				14'b11101011001111: Data_out <= 16'hC18E	;
				14'b11101011010000: Data_out <= 16'hC199	;
				14'b11101011010001: Data_out <= 16'hC1A4	;
				14'b11101011010010: Data_out <= 16'hC1AE	;
				14'b11101011010011: Data_out <= 16'hC1B9	;
				14'b11101011010100: Data_out <= 16'hC1C4	;
				14'b11101011010101: Data_out <= 16'hC1CF	;
				14'b11101011010110: Data_out <= 16'hC1DA	;
				14'b11101011010111: Data_out <= 16'hC1E5	;
				14'b11101011011000: Data_out <= 16'hC1F0	;
				14'b11101011011001: Data_out <= 16'hC1FB	;
				14'b11101011011010: Data_out <= 16'hC206	;
				14'b11101011011011: Data_out <= 16'hC211	;
				14'b11101011011100: Data_out <= 16'hC21C	;
				14'b11101011011101: Data_out <= 16'hC227	;
				14'b11101011011110: Data_out <= 16'hC232	;
				14'b11101011011111: Data_out <= 16'hC23D	;
				14'b11101011100000: Data_out <= 16'hC248	;
				14'b11101011100001: Data_out <= 16'hC253	;
				14'b11101011100010: Data_out <= 16'hC25E	;
				14'b11101011100011: Data_out <= 16'hC269	;
				14'b11101011100100: Data_out <= 16'hC274	;
				14'b11101011100101: Data_out <= 16'hC27F	;
				14'b11101011100110: Data_out <= 16'hC28A	;
				14'b11101011100111: Data_out <= 16'hC296	;
				14'b11101011101000: Data_out <= 16'hC2A1	;
				14'b11101011101001: Data_out <= 16'hC2AC	;
				14'b11101011101010: Data_out <= 16'hC2B7	;
				14'b11101011101011: Data_out <= 16'hC2C2	;
				14'b11101011101100: Data_out <= 16'hC2CD	;
				14'b11101011101101: Data_out <= 16'hC2D8	;
				14'b11101011101110: Data_out <= 16'hC2E3	;
				14'b11101011101111: Data_out <= 16'hC2EE	;
				14'b11101011110000: Data_out <= 16'hC2F9	;
				14'b11101011110001: Data_out <= 16'hC304	;
				14'b11101011110010: Data_out <= 16'hC30F	;
				14'b11101011110011: Data_out <= 16'hC31A	;
				14'b11101011110100: Data_out <= 16'hC325	;
				14'b11101011110101: Data_out <= 16'hC330	;
				14'b11101011110110: Data_out <= 16'hC33B	;
				14'b11101011110111: Data_out <= 16'hC346	;
				14'b11101011111000: Data_out <= 16'hC351	;
				14'b11101011111001: Data_out <= 16'hC35C	;
				14'b11101011111010: Data_out <= 16'hC367	;
				14'b11101011111011: Data_out <= 16'hC372	;
				14'b11101011111100: Data_out <= 16'hC37E	;
				14'b11101011111101: Data_out <= 16'hC389	;
				14'b11101011111110: Data_out <= 16'hC394	;
				14'b11101011111111: Data_out <= 16'hC39F	;
				14'b11101100000000: Data_out <= 16'hC3AA	;
				14'b11101100000001: Data_out <= 16'hC3B5	;
				14'b11101100000010: Data_out <= 16'hC3C0	;
				14'b11101100000011: Data_out <= 16'hC3CB	;
				14'b11101100000100: Data_out <= 16'hC3D6	;
				14'b11101100000101: Data_out <= 16'hC3E1	;
				14'b11101100000110: Data_out <= 16'hC3EC	;
				14'b11101100000111: Data_out <= 16'hC3F7	;
				14'b11101100001000: Data_out <= 16'hC403	;
				14'b11101100001001: Data_out <= 16'hC40E	;
				14'b11101100001010: Data_out <= 16'hC419	;
				14'b11101100001011: Data_out <= 16'hC424	;
				14'b11101100001100: Data_out <= 16'hC42F	;
				14'b11101100001101: Data_out <= 16'hC43A	;
				14'b11101100001110: Data_out <= 16'hC445	;
				14'b11101100001111: Data_out <= 16'hC450	;
				14'b11101100010000: Data_out <= 16'hC45B	;
				14'b11101100010001: Data_out <= 16'hC467	;
				14'b11101100010010: Data_out <= 16'hC472	;
				14'b11101100010011: Data_out <= 16'hC47D	;
				14'b11101100010100: Data_out <= 16'hC488	;
				14'b11101100010101: Data_out <= 16'hC493	;
				14'b11101100010110: Data_out <= 16'hC49E	;
				14'b11101100010111: Data_out <= 16'hC4A9	;
				14'b11101100011000: Data_out <= 16'hC4B4	;
				14'b11101100011001: Data_out <= 16'hC4C0	;
				14'b11101100011010: Data_out <= 16'hC4CB	;
				14'b11101100011011: Data_out <= 16'hC4D6	;
				14'b11101100011100: Data_out <= 16'hC4E1	;
				14'b11101100011101: Data_out <= 16'hC4EC	;
				14'b11101100011110: Data_out <= 16'hC4F7	;
				14'b11101100011111: Data_out <= 16'hC502	;
				14'b11101100100000: Data_out <= 16'hC50E	;
				14'b11101100100001: Data_out <= 16'hC519	;
				14'b11101100100010: Data_out <= 16'hC524	;
				14'b11101100100011: Data_out <= 16'hC52F	;
				14'b11101100100100: Data_out <= 16'hC53A	;
				14'b11101100100101: Data_out <= 16'hC545	;
				14'b11101100100110: Data_out <= 16'hC551	;
				14'b11101100100111: Data_out <= 16'hC55C	;
				14'b11101100101000: Data_out <= 16'hC567	;
				14'b11101100101001: Data_out <= 16'hC572	;
				14'b11101100101010: Data_out <= 16'hC57D	;
				14'b11101100101011: Data_out <= 16'hC588	;
				14'b11101100101100: Data_out <= 16'hC594	;
				14'b11101100101101: Data_out <= 16'hC59F	;
				14'b11101100101110: Data_out <= 16'hC5AA	;
				14'b11101100101111: Data_out <= 16'hC5B5	;
				14'b11101100110000: Data_out <= 16'hC5C0	;
				14'b11101100110001: Data_out <= 16'hC5CC	;
				14'b11101100110010: Data_out <= 16'hC5D7	;
				14'b11101100110011: Data_out <= 16'hC5E2	;
				14'b11101100110100: Data_out <= 16'hC5ED	;
				14'b11101100110101: Data_out <= 16'hC5F8	;
				14'b11101100110110: Data_out <= 16'hC604	;
				14'b11101100110111: Data_out <= 16'hC60F	;
				14'b11101100111000: Data_out <= 16'hC61A	;
				14'b11101100111001: Data_out <= 16'hC625	;
				14'b11101100111010: Data_out <= 16'hC630	;
				14'b11101100111011: Data_out <= 16'hC63C	;
				14'b11101100111100: Data_out <= 16'hC647	;
				14'b11101100111101: Data_out <= 16'hC652	;
				14'b11101100111110: Data_out <= 16'hC65D	;
				14'b11101100111111: Data_out <= 16'hC668	;
				14'b11101101000000: Data_out <= 16'hC674	;
				14'b11101101000001: Data_out <= 16'hC67F	;
				14'b11101101000010: Data_out <= 16'hC68A	;
				14'b11101101000011: Data_out <= 16'hC695	;
				14'b11101101000100: Data_out <= 16'hC6A1	;
				14'b11101101000101: Data_out <= 16'hC6AC	;
				14'b11101101000110: Data_out <= 16'hC6B7	;
				14'b11101101000111: Data_out <= 16'hC6C2	;
				14'b11101101001000: Data_out <= 16'hC6CE	;
				14'b11101101001001: Data_out <= 16'hC6D9	;
				14'b11101101001010: Data_out <= 16'hC6E4	;
				14'b11101101001011: Data_out <= 16'hC6EF	;
				14'b11101101001100: Data_out <= 16'hC6FB	;
				14'b11101101001101: Data_out <= 16'hC706	;
				14'b11101101001110: Data_out <= 16'hC711	;
				14'b11101101001111: Data_out <= 16'hC71C	;
				14'b11101101010000: Data_out <= 16'hC728	;
				14'b11101101010001: Data_out <= 16'hC733	;
				14'b11101101010010: Data_out <= 16'hC73E	;
				14'b11101101010011: Data_out <= 16'hC749	;
				14'b11101101010100: Data_out <= 16'hC755	;
				14'b11101101010101: Data_out <= 16'hC760	;
				14'b11101101010110: Data_out <= 16'hC76B	;
				14'b11101101010111: Data_out <= 16'hC776	;
				14'b11101101011000: Data_out <= 16'hC782	;
				14'b11101101011001: Data_out <= 16'hC78D	;
				14'b11101101011010: Data_out <= 16'hC798	;
				14'b11101101011011: Data_out <= 16'hC7A4	;
				14'b11101101011100: Data_out <= 16'hC7AF	;
				14'b11101101011101: Data_out <= 16'hC7BA	;
				14'b11101101011110: Data_out <= 16'hC7C5	;
				14'b11101101011111: Data_out <= 16'hC7D1	;
				14'b11101101100000: Data_out <= 16'hC7DC	;
				14'b11101101100001: Data_out <= 16'hC7E7	;
				14'b11101101100010: Data_out <= 16'hC7F3	;
				14'b11101101100011: Data_out <= 16'hC7FE	;
				14'b11101101100100: Data_out <= 16'hC809	;
				14'b11101101100101: Data_out <= 16'hC814	;
				14'b11101101100110: Data_out <= 16'hC820	;
				14'b11101101100111: Data_out <= 16'hC82B	;
				14'b11101101101000: Data_out <= 16'hC836	;
				14'b11101101101001: Data_out <= 16'hC842	;
				14'b11101101101010: Data_out <= 16'hC84D	;
				14'b11101101101011: Data_out <= 16'hC858	;
				14'b11101101101100: Data_out <= 16'hC864	;
				14'b11101101101101: Data_out <= 16'hC86F	;
				14'b11101101101110: Data_out <= 16'hC87A	;
				14'b11101101101111: Data_out <= 16'hC886	;
				14'b11101101110000: Data_out <= 16'hC891	;
				14'b11101101110001: Data_out <= 16'hC89C	;
				14'b11101101110010: Data_out <= 16'hC8A8	;
				14'b11101101110011: Data_out <= 16'hC8B3	;
				14'b11101101110100: Data_out <= 16'hC8BE	;
				14'b11101101110101: Data_out <= 16'hC8CA	;
				14'b11101101110110: Data_out <= 16'hC8D5	;
				14'b11101101110111: Data_out <= 16'hC8E0	;
				14'b11101101111000: Data_out <= 16'hC8EC	;
				14'b11101101111001: Data_out <= 16'hC8F7	;
				14'b11101101111010: Data_out <= 16'hC902	;
				14'b11101101111011: Data_out <= 16'hC90E	;
				14'b11101101111100: Data_out <= 16'hC919	;
				14'b11101101111101: Data_out <= 16'hC924	;
				14'b11101101111110: Data_out <= 16'hC930	;
				14'b11101101111111: Data_out <= 16'hC93B	;
				14'b11101110000000: Data_out <= 16'hC946	;
				14'b11101110000001: Data_out <= 16'hC952	;
				14'b11101110000010: Data_out <= 16'hC95D	;
				14'b11101110000011: Data_out <= 16'hC968	;
				14'b11101110000100: Data_out <= 16'hC974	;
				14'b11101110000101: Data_out <= 16'hC97F	;
				14'b11101110000110: Data_out <= 16'hC98B	;
				14'b11101110000111: Data_out <= 16'hC996	;
				14'b11101110001000: Data_out <= 16'hC9A1	;
				14'b11101110001001: Data_out <= 16'hC9AD	;
				14'b11101110001010: Data_out <= 16'hC9B8	;
				14'b11101110001011: Data_out <= 16'hC9C3	;
				14'b11101110001100: Data_out <= 16'hC9CF	;
				14'b11101110001101: Data_out <= 16'hC9DA	;
				14'b11101110001110: Data_out <= 16'hC9E6	;
				14'b11101110001111: Data_out <= 16'hC9F1	;
				14'b11101110010000: Data_out <= 16'hC9FC	;
				14'b11101110010001: Data_out <= 16'hCA08	;
				14'b11101110010010: Data_out <= 16'hCA13	;
				14'b11101110010011: Data_out <= 16'hCA1F	;
				14'b11101110010100: Data_out <= 16'hCA2A	;
				14'b11101110010101: Data_out <= 16'hCA35	;
				14'b11101110010110: Data_out <= 16'hCA41	;
				14'b11101110010111: Data_out <= 16'hCA4C	;
				14'b11101110011000: Data_out <= 16'hCA58	;
				14'b11101110011001: Data_out <= 16'hCA63	;
				14'b11101110011010: Data_out <= 16'hCA6E	;
				14'b11101110011011: Data_out <= 16'hCA7A	;
				14'b11101110011100: Data_out <= 16'hCA85	;
				14'b11101110011101: Data_out <= 16'hCA91	;
				14'b11101110011110: Data_out <= 16'hCA9C	;
				14'b11101110011111: Data_out <= 16'hCAA8	;
				14'b11101110100000: Data_out <= 16'hCAB3	;
				14'b11101110100001: Data_out <= 16'hCABE	;
				14'b11101110100010: Data_out <= 16'hCACA	;
				14'b11101110100011: Data_out <= 16'hCAD5	;
				14'b11101110100100: Data_out <= 16'hCAE1	;
				14'b11101110100101: Data_out <= 16'hCAEC	;
				14'b11101110100110: Data_out <= 16'hCAF8	;
				14'b11101110100111: Data_out <= 16'hCB03	;
				14'b11101110101000: Data_out <= 16'hCB0E	;
				14'b11101110101001: Data_out <= 16'hCB1A	;
				14'b11101110101010: Data_out <= 16'hCB25	;
				14'b11101110101011: Data_out <= 16'hCB31	;
				14'b11101110101100: Data_out <= 16'hCB3C	;
				14'b11101110101101: Data_out <= 16'hCB48	;
				14'b11101110101110: Data_out <= 16'hCB53	;
				14'b11101110101111: Data_out <= 16'hCB5F	;
				14'b11101110110000: Data_out <= 16'hCB6A	;
				14'b11101110110001: Data_out <= 16'hCB75	;
				14'b11101110110010: Data_out <= 16'hCB81	;
				14'b11101110110011: Data_out <= 16'hCB8C	;
				14'b11101110110100: Data_out <= 16'hCB98	;
				14'b11101110110101: Data_out <= 16'hCBA3	;
				14'b11101110110110: Data_out <= 16'hCBAF	;
				14'b11101110110111: Data_out <= 16'hCBBA	;
				14'b11101110111000: Data_out <= 16'hCBC6	;
				14'b11101110111001: Data_out <= 16'hCBD1	;
				14'b11101110111010: Data_out <= 16'hCBDD	;
				14'b11101110111011: Data_out <= 16'hCBE8	;
				14'b11101110111100: Data_out <= 16'hCBF4	;
				14'b11101110111101: Data_out <= 16'hCBFF	;
				14'b11101110111110: Data_out <= 16'hCC0B	;
				14'b11101110111111: Data_out <= 16'hCC16	;
				14'b11101111000000: Data_out <= 16'hCC22	;
				14'b11101111000001: Data_out <= 16'hCC2D	;
				14'b11101111000010: Data_out <= 16'hCC39	;
				14'b11101111000011: Data_out <= 16'hCC44	;
				14'b11101111000100: Data_out <= 16'hCC50	;
				14'b11101111000101: Data_out <= 16'hCC5B	;
				14'b11101111000110: Data_out <= 16'hCC67	;
				14'b11101111000111: Data_out <= 16'hCC72	;
				14'b11101111001000: Data_out <= 16'hCC7E	;
				14'b11101111001001: Data_out <= 16'hCC89	;
				14'b11101111001010: Data_out <= 16'hCC95	;
				14'b11101111001011: Data_out <= 16'hCCA0	;
				14'b11101111001100: Data_out <= 16'hCCAC	;
				14'b11101111001101: Data_out <= 16'hCCB7	;
				14'b11101111001110: Data_out <= 16'hCCC3	;
				14'b11101111001111: Data_out <= 16'hCCCE	;
				14'b11101111010000: Data_out <= 16'hCCDA	;
				14'b11101111010001: Data_out <= 16'hCCE5	;
				14'b11101111010010: Data_out <= 16'hCCF1	;
				14'b11101111010011: Data_out <= 16'hCCFC	;
				14'b11101111010100: Data_out <= 16'hCD08	;
				14'b11101111010101: Data_out <= 16'hCD13	;
				14'b11101111010110: Data_out <= 16'hCD1F	;
				14'b11101111010111: Data_out <= 16'hCD2A	;
				14'b11101111011000: Data_out <= 16'hCD36	;
				14'b11101111011001: Data_out <= 16'hCD41	;
				14'b11101111011010: Data_out <= 16'hCD4D	;
				14'b11101111011011: Data_out <= 16'hCD58	;
				14'b11101111011100: Data_out <= 16'hCD64	;
				14'b11101111011101: Data_out <= 16'hCD70	;
				14'b11101111011110: Data_out <= 16'hCD7B	;
				14'b11101111011111: Data_out <= 16'hCD87	;
				14'b11101111100000: Data_out <= 16'hCD92	;
				14'b11101111100001: Data_out <= 16'hCD9E	;
				14'b11101111100010: Data_out <= 16'hCDA9	;
				14'b11101111100011: Data_out <= 16'hCDB5	;
				14'b11101111100100: Data_out <= 16'hCDC0	;
				14'b11101111100101: Data_out <= 16'hCDCC	;
				14'b11101111100110: Data_out <= 16'hCDD7	;
				14'b11101111100111: Data_out <= 16'hCDE3	;
				14'b11101111101000: Data_out <= 16'hCDEF	;
				14'b11101111101001: Data_out <= 16'hCDFA	;
				14'b11101111101010: Data_out <= 16'hCE06	;
				14'b11101111101011: Data_out <= 16'hCE11	;
				14'b11101111101100: Data_out <= 16'hCE1D	;
				14'b11101111101101: Data_out <= 16'hCE28	;
				14'b11101111101110: Data_out <= 16'hCE34	;
				14'b11101111101111: Data_out <= 16'hCE40	;
				14'b11101111110000: Data_out <= 16'hCE4B	;
				14'b11101111110001: Data_out <= 16'hCE57	;
				14'b11101111110010: Data_out <= 16'hCE62	;
				14'b11101111110011: Data_out <= 16'hCE6E	;
				14'b11101111110100: Data_out <= 16'hCE7A	;
				14'b11101111110101: Data_out <= 16'hCE85	;
				14'b11101111110110: Data_out <= 16'hCE91	;
				14'b11101111110111: Data_out <= 16'hCE9C	;
				14'b11101111111000: Data_out <= 16'hCEA8	;
				14'b11101111111001: Data_out <= 16'hCEB3	;
				14'b11101111111010: Data_out <= 16'hCEBF	;
				14'b11101111111011: Data_out <= 16'hCECB	;
				14'b11101111111100: Data_out <= 16'hCED6	;
				14'b11101111111101: Data_out <= 16'hCEE2	;
				14'b11101111111110: Data_out <= 16'hCEED	;
				14'b11101111111111: Data_out <= 16'hCEF9	;
				14'b11110000000000: Data_out <= 16'hCF05	;
				14'b11110000000001: Data_out <= 16'hCF10	;
				14'b11110000000010: Data_out <= 16'hCF1C	;
				14'b11110000000011: Data_out <= 16'hCF28	;
				14'b11110000000100: Data_out <= 16'hCF33	;
				14'b11110000000101: Data_out <= 16'hCF3F	;
				14'b11110000000110: Data_out <= 16'hCF4A	;
				14'b11110000000111: Data_out <= 16'hCF56	;
				14'b11110000001000: Data_out <= 16'hCF62	;
				14'b11110000001001: Data_out <= 16'hCF6D	;
				14'b11110000001010: Data_out <= 16'hCF79	;
				14'b11110000001011: Data_out <= 16'hCF85	;
				14'b11110000001100: Data_out <= 16'hCF90	;
				14'b11110000001101: Data_out <= 16'hCF9C	;
				14'b11110000001110: Data_out <= 16'hCFA7	;
				14'b11110000001111: Data_out <= 16'hCFB3	;
				14'b11110000010000: Data_out <= 16'hCFBF	;
				14'b11110000010001: Data_out <= 16'hCFCA	;
				14'b11110000010010: Data_out <= 16'hCFD6	;
				14'b11110000010011: Data_out <= 16'hCFE2	;
				14'b11110000010100: Data_out <= 16'hCFED	;
				14'b11110000010101: Data_out <= 16'hCFF9	;
				14'b11110000010110: Data_out <= 16'hD005	;
				14'b11110000010111: Data_out <= 16'hD010	;
				14'b11110000011000: Data_out <= 16'hD01C	;
				14'b11110000011001: Data_out <= 16'hD028	;
				14'b11110000011010: Data_out <= 16'hD033	;
				14'b11110000011011: Data_out <= 16'hD03F	;
				14'b11110000011100: Data_out <= 16'hD04A	;
				14'b11110000011101: Data_out <= 16'hD056	;
				14'b11110000011110: Data_out <= 16'hD062	;
				14'b11110000011111: Data_out <= 16'hD06D	;
				14'b11110000100000: Data_out <= 16'hD079	;
				14'b11110000100001: Data_out <= 16'hD085	;
				14'b11110000100010: Data_out <= 16'hD090	;
				14'b11110000100011: Data_out <= 16'hD09C	;
				14'b11110000100100: Data_out <= 16'hD0A8	;
				14'b11110000100101: Data_out <= 16'hD0B4	;
				14'b11110000100110: Data_out <= 16'hD0BF	;
				14'b11110000100111: Data_out <= 16'hD0CB	;
				14'b11110000101000: Data_out <= 16'hD0D7	;
				14'b11110000101001: Data_out <= 16'hD0E2	;
				14'b11110000101010: Data_out <= 16'hD0EE	;
				14'b11110000101011: Data_out <= 16'hD0FA	;
				14'b11110000101100: Data_out <= 16'hD105	;
				14'b11110000101101: Data_out <= 16'hD111	;
				14'b11110000101110: Data_out <= 16'hD11D	;
				14'b11110000101111: Data_out <= 16'hD128	;
				14'b11110000110000: Data_out <= 16'hD134	;
				14'b11110000110001: Data_out <= 16'hD140	;
				14'b11110000110010: Data_out <= 16'hD14B	;
				14'b11110000110011: Data_out <= 16'hD157	;
				14'b11110000110100: Data_out <= 16'hD163	;
				14'b11110000110101: Data_out <= 16'hD16F	;
				14'b11110000110110: Data_out <= 16'hD17A	;
				14'b11110000110111: Data_out <= 16'hD186	;
				14'b11110000111000: Data_out <= 16'hD192	;
				14'b11110000111001: Data_out <= 16'hD19D	;
				14'b11110000111010: Data_out <= 16'hD1A9	;
				14'b11110000111011: Data_out <= 16'hD1B5	;
				14'b11110000111100: Data_out <= 16'hD1C1	;
				14'b11110000111101: Data_out <= 16'hD1CC	;
				14'b11110000111110: Data_out <= 16'hD1D8	;
				14'b11110000111111: Data_out <= 16'hD1E4	;
				14'b11110001000000: Data_out <= 16'hD1EF	;
				14'b11110001000001: Data_out <= 16'hD1FB	;
				14'b11110001000010: Data_out <= 16'hD207	;
				14'b11110001000011: Data_out <= 16'hD213	;
				14'b11110001000100: Data_out <= 16'hD21E	;
				14'b11110001000101: Data_out <= 16'hD22A	;
				14'b11110001000110: Data_out <= 16'hD236	;
				14'b11110001000111: Data_out <= 16'hD242	;
				14'b11110001001000: Data_out <= 16'hD24D	;
				14'b11110001001001: Data_out <= 16'hD259	;
				14'b11110001001010: Data_out <= 16'hD265	;
				14'b11110001001011: Data_out <= 16'hD270	;
				14'b11110001001100: Data_out <= 16'hD27C	;
				14'b11110001001101: Data_out <= 16'hD288	;
				14'b11110001001110: Data_out <= 16'hD294	;
				14'b11110001001111: Data_out <= 16'hD29F	;
				14'b11110001010000: Data_out <= 16'hD2AB	;
				14'b11110001010001: Data_out <= 16'hD2B7	;
				14'b11110001010010: Data_out <= 16'hD2C3	;
				14'b11110001010011: Data_out <= 16'hD2CE	;
				14'b11110001010100: Data_out <= 16'hD2DA	;
				14'b11110001010101: Data_out <= 16'hD2E6	;
				14'b11110001010110: Data_out <= 16'hD2F2	;
				14'b11110001010111: Data_out <= 16'hD2FE	;
				14'b11110001011000: Data_out <= 16'hD309	;
				14'b11110001011001: Data_out <= 16'hD315	;
				14'b11110001011010: Data_out <= 16'hD321	;
				14'b11110001011011: Data_out <= 16'hD32D	;
				14'b11110001011100: Data_out <= 16'hD338	;
				14'b11110001011101: Data_out <= 16'hD344	;
				14'b11110001011110: Data_out <= 16'hD350	;
				14'b11110001011111: Data_out <= 16'hD35C	;
				14'b11110001100000: Data_out <= 16'hD367	;
				14'b11110001100001: Data_out <= 16'hD373	;
				14'b11110001100010: Data_out <= 16'hD37F	;
				14'b11110001100011: Data_out <= 16'hD38B	;
				14'b11110001100100: Data_out <= 16'hD397	;
				14'b11110001100101: Data_out <= 16'hD3A2	;
				14'b11110001100110: Data_out <= 16'hD3AE	;
				14'b11110001100111: Data_out <= 16'hD3BA	;
				14'b11110001101000: Data_out <= 16'hD3C6	;
				14'b11110001101001: Data_out <= 16'hD3D2	;
				14'b11110001101010: Data_out <= 16'hD3DD	;
				14'b11110001101011: Data_out <= 16'hD3E9	;
				14'b11110001101100: Data_out <= 16'hD3F5	;
				14'b11110001101101: Data_out <= 16'hD401	;
				14'b11110001101110: Data_out <= 16'hD40D	;
				14'b11110001101111: Data_out <= 16'hD418	;
				14'b11110001110000: Data_out <= 16'hD424	;
				14'b11110001110001: Data_out <= 16'hD430	;
				14'b11110001110010: Data_out <= 16'hD43C	;
				14'b11110001110011: Data_out <= 16'hD448	;
				14'b11110001110100: Data_out <= 16'hD453	;
				14'b11110001110101: Data_out <= 16'hD45F	;
				14'b11110001110110: Data_out <= 16'hD46B	;
				14'b11110001110111: Data_out <= 16'hD477	;
				14'b11110001111000: Data_out <= 16'hD483	;
				14'b11110001111001: Data_out <= 16'hD48E	;
				14'b11110001111010: Data_out <= 16'hD49A	;
				14'b11110001111011: Data_out <= 16'hD4A6	;
				14'b11110001111100: Data_out <= 16'hD4B2	;
				14'b11110001111101: Data_out <= 16'hD4BE	;
				14'b11110001111110: Data_out <= 16'hD4CA	;
				14'b11110001111111: Data_out <= 16'hD4D5	;
				14'b11110010000000: Data_out <= 16'hD4E1	;
				14'b11110010000001: Data_out <= 16'hD4ED	;
				14'b11110010000010: Data_out <= 16'hD4F9	;
				14'b11110010000011: Data_out <= 16'hD505	;
				14'b11110010000100: Data_out <= 16'hD511	;
				14'b11110010000101: Data_out <= 16'hD51C	;
				14'b11110010000110: Data_out <= 16'hD528	;
				14'b11110010000111: Data_out <= 16'hD534	;
				14'b11110010001000: Data_out <= 16'hD540	;
				14'b11110010001001: Data_out <= 16'hD54C	;
				14'b11110010001010: Data_out <= 16'hD558	;
				14'b11110010001011: Data_out <= 16'hD563	;
				14'b11110010001100: Data_out <= 16'hD56F	;
				14'b11110010001101: Data_out <= 16'hD57B	;
				14'b11110010001110: Data_out <= 16'hD587	;
				14'b11110010001111: Data_out <= 16'hD593	;
				14'b11110010010000: Data_out <= 16'hD59F	;
				14'b11110010010001: Data_out <= 16'hD5AB	;
				14'b11110010010010: Data_out <= 16'hD5B6	;
				14'b11110010010011: Data_out <= 16'hD5C2	;
				14'b11110010010100: Data_out <= 16'hD5CE	;
				14'b11110010010101: Data_out <= 16'hD5DA	;
				14'b11110010010110: Data_out <= 16'hD5E6	;
				14'b11110010010111: Data_out <= 16'hD5F2	;
				14'b11110010011000: Data_out <= 16'hD5FE	;
				14'b11110010011001: Data_out <= 16'hD60A	;
				14'b11110010011010: Data_out <= 16'hD615	;
				14'b11110010011011: Data_out <= 16'hD621	;
				14'b11110010011100: Data_out <= 16'hD62D	;
				14'b11110010011101: Data_out <= 16'hD639	;
				14'b11110010011110: Data_out <= 16'hD645	;
				14'b11110010011111: Data_out <= 16'hD651	;
				14'b11110010100000: Data_out <= 16'hD65D	;
				14'b11110010100001: Data_out <= 16'hD669	;
				14'b11110010100010: Data_out <= 16'hD674	;
				14'b11110010100011: Data_out <= 16'hD680	;
				14'b11110010100100: Data_out <= 16'hD68C	;
				14'b11110010100101: Data_out <= 16'hD698	;
				14'b11110010100110: Data_out <= 16'hD6A4	;
				14'b11110010100111: Data_out <= 16'hD6B0	;
				14'b11110010101000: Data_out <= 16'hD6BC	;
				14'b11110010101001: Data_out <= 16'hD6C8	;
				14'b11110010101010: Data_out <= 16'hD6D4	;
				14'b11110010101011: Data_out <= 16'hD6DF	;
				14'b11110010101100: Data_out <= 16'hD6EB	;
				14'b11110010101101: Data_out <= 16'hD6F7	;
				14'b11110010101110: Data_out <= 16'hD703	;
				14'b11110010101111: Data_out <= 16'hD70F	;
				14'b11110010110000: Data_out <= 16'hD71B	;
				14'b11110010110001: Data_out <= 16'hD727	;
				14'b11110010110010: Data_out <= 16'hD733	;
				14'b11110010110011: Data_out <= 16'hD73F	;
				14'b11110010110100: Data_out <= 16'hD74B	;
				14'b11110010110101: Data_out <= 16'hD757	;
				14'b11110010110110: Data_out <= 16'hD762	;
				14'b11110010110111: Data_out <= 16'hD76E	;
				14'b11110010111000: Data_out <= 16'hD77A	;
				14'b11110010111001: Data_out <= 16'hD786	;
				14'b11110010111010: Data_out <= 16'hD792	;
				14'b11110010111011: Data_out <= 16'hD79E	;
				14'b11110010111100: Data_out <= 16'hD7AA	;
				14'b11110010111101: Data_out <= 16'hD7B6	;
				14'b11110010111110: Data_out <= 16'hD7C2	;
				14'b11110010111111: Data_out <= 16'hD7CE	;
				14'b11110011000000: Data_out <= 16'hD7DA	;
				14'b11110011000001: Data_out <= 16'hD7E6	;
				14'b11110011000010: Data_out <= 16'hD7F2	;
				14'b11110011000011: Data_out <= 16'hD7FD	;
				14'b11110011000100: Data_out <= 16'hD809	;
				14'b11110011000101: Data_out <= 16'hD815	;
				14'b11110011000110: Data_out <= 16'hD821	;
				14'b11110011000111: Data_out <= 16'hD82D	;
				14'b11110011001000: Data_out <= 16'hD839	;
				14'b11110011001001: Data_out <= 16'hD845	;
				14'b11110011001010: Data_out <= 16'hD851	;
				14'b11110011001011: Data_out <= 16'hD85D	;
				14'b11110011001100: Data_out <= 16'hD869	;
				14'b11110011001101: Data_out <= 16'hD875	;
				14'b11110011001110: Data_out <= 16'hD881	;
				14'b11110011001111: Data_out <= 16'hD88D	;
				14'b11110011010000: Data_out <= 16'hD899	;
				14'b11110011010001: Data_out <= 16'hD8A5	;
				14'b11110011010010: Data_out <= 16'hD8B1	;
				14'b11110011010011: Data_out <= 16'hD8BD	;
				14'b11110011010100: Data_out <= 16'hD8C9	;
				14'b11110011010101: Data_out <= 16'hD8D5	;
				14'b11110011010110: Data_out <= 16'hD8E1	;
				14'b11110011010111: Data_out <= 16'hD8ED	;
				14'b11110011011000: Data_out <= 16'hD8F8	;
				14'b11110011011001: Data_out <= 16'hD904	;
				14'b11110011011010: Data_out <= 16'hD910	;
				14'b11110011011011: Data_out <= 16'hD91C	;
				14'b11110011011100: Data_out <= 16'hD928	;
				14'b11110011011101: Data_out <= 16'hD934	;
				14'b11110011011110: Data_out <= 16'hD940	;
				14'b11110011011111: Data_out <= 16'hD94C	;
				14'b11110011100000: Data_out <= 16'hD958	;
				14'b11110011100001: Data_out <= 16'hD964	;
				14'b11110011100010: Data_out <= 16'hD970	;
				14'b11110011100011: Data_out <= 16'hD97C	;
				14'b11110011100100: Data_out <= 16'hD988	;
				14'b11110011100101: Data_out <= 16'hD994	;
				14'b11110011100110: Data_out <= 16'hD9A0	;
				14'b11110011100111: Data_out <= 16'hD9AC	;
				14'b11110011101000: Data_out <= 16'hD9B8	;
				14'b11110011101001: Data_out <= 16'hD9C4	;
				14'b11110011101010: Data_out <= 16'hD9D0	;
				14'b11110011101011: Data_out <= 16'hD9DC	;
				14'b11110011101100: Data_out <= 16'hD9E8	;
				14'b11110011101101: Data_out <= 16'hD9F4	;
				14'b11110011101110: Data_out <= 16'hDA00	;
				14'b11110011101111: Data_out <= 16'hDA0C	;
				14'b11110011110000: Data_out <= 16'hDA18	;
				14'b11110011110001: Data_out <= 16'hDA24	;
				14'b11110011110010: Data_out <= 16'hDA30	;
				14'b11110011110011: Data_out <= 16'hDA3C	;
				14'b11110011110100: Data_out <= 16'hDA48	;
				14'b11110011110101: Data_out <= 16'hDA54	;
				14'b11110011110110: Data_out <= 16'hDA60	;
				14'b11110011110111: Data_out <= 16'hDA6C	;
				14'b11110011111000: Data_out <= 16'hDA78	;
				14'b11110011111001: Data_out <= 16'hDA84	;
				14'b11110011111010: Data_out <= 16'hDA90	;
				14'b11110011111011: Data_out <= 16'hDA9C	;
				14'b11110011111100: Data_out <= 16'hDAA8	;
				14'b11110011111101: Data_out <= 16'hDAB4	;
				14'b11110011111110: Data_out <= 16'hDAC0	;
				14'b11110011111111: Data_out <= 16'hDACC	;
				14'b11110100000000: Data_out <= 16'hDAD8	;
				14'b11110100000001: Data_out <= 16'hDAE4	;
				14'b11110100000010: Data_out <= 16'hDAF0	;
				14'b11110100000011: Data_out <= 16'hDAFC	;
				14'b11110100000100: Data_out <= 16'hDB08	;
				14'b11110100000101: Data_out <= 16'hDB14	;
				14'b11110100000110: Data_out <= 16'hDB21	;
				14'b11110100000111: Data_out <= 16'hDB2D	;
				14'b11110100001000: Data_out <= 16'hDB39	;
				14'b11110100001001: Data_out <= 16'hDB45	;
				14'b11110100001010: Data_out <= 16'hDB51	;
				14'b11110100001011: Data_out <= 16'hDB5D	;
				14'b11110100001100: Data_out <= 16'hDB69	;
				14'b11110100001101: Data_out <= 16'hDB75	;
				14'b11110100001110: Data_out <= 16'hDB81	;
				14'b11110100001111: Data_out <= 16'hDB8D	;
				14'b11110100010000: Data_out <= 16'hDB99	;
				14'b11110100010001: Data_out <= 16'hDBA5	;
				14'b11110100010010: Data_out <= 16'hDBB1	;
				14'b11110100010011: Data_out <= 16'hDBBD	;
				14'b11110100010100: Data_out <= 16'hDBC9	;
				14'b11110100010101: Data_out <= 16'hDBD5	;
				14'b11110100010110: Data_out <= 16'hDBE1	;
				14'b11110100010111: Data_out <= 16'hDBED	;
				14'b11110100011000: Data_out <= 16'hDBF9	;
				14'b11110100011001: Data_out <= 16'hDC05	;
				14'b11110100011010: Data_out <= 16'hDC11	;
				14'b11110100011011: Data_out <= 16'hDC1E	;
				14'b11110100011100: Data_out <= 16'hDC2A	;
				14'b11110100011101: Data_out <= 16'hDC36	;
				14'b11110100011110: Data_out <= 16'hDC42	;
				14'b11110100011111: Data_out <= 16'hDC4E	;
				14'b11110100100000: Data_out <= 16'hDC5A	;
				14'b11110100100001: Data_out <= 16'hDC66	;
				14'b11110100100010: Data_out <= 16'hDC72	;
				14'b11110100100011: Data_out <= 16'hDC7E	;
				14'b11110100100100: Data_out <= 16'hDC8A	;
				14'b11110100100101: Data_out <= 16'hDC96	;
				14'b11110100100110: Data_out <= 16'hDCA2	;
				14'b11110100100111: Data_out <= 16'hDCAE	;
				14'b11110100101000: Data_out <= 16'hDCBA	;
				14'b11110100101001: Data_out <= 16'hDCC7	;
				14'b11110100101010: Data_out <= 16'hDCD3	;
				14'b11110100101011: Data_out <= 16'hDCDF	;
				14'b11110100101100: Data_out <= 16'hDCEB	;
				14'b11110100101101: Data_out <= 16'hDCF7	;
				14'b11110100101110: Data_out <= 16'hDD03	;
				14'b11110100101111: Data_out <= 16'hDD0F	;
				14'b11110100110000: Data_out <= 16'hDD1B	;
				14'b11110100110001: Data_out <= 16'hDD27	;
				14'b11110100110010: Data_out <= 16'hDD33	;
				14'b11110100110011: Data_out <= 16'hDD3F	;
				14'b11110100110100: Data_out <= 16'hDD4B	;
				14'b11110100110101: Data_out <= 16'hDD58	;
				14'b11110100110110: Data_out <= 16'hDD64	;
				14'b11110100110111: Data_out <= 16'hDD70	;
				14'b11110100111000: Data_out <= 16'hDD7C	;
				14'b11110100111001: Data_out <= 16'hDD88	;
				14'b11110100111010: Data_out <= 16'hDD94	;
				14'b11110100111011: Data_out <= 16'hDDA0	;
				14'b11110100111100: Data_out <= 16'hDDAC	;
				14'b11110100111101: Data_out <= 16'hDDB8	;
				14'b11110100111110: Data_out <= 16'hDDC5	;
				14'b11110100111111: Data_out <= 16'hDDD1	;
				14'b11110101000000: Data_out <= 16'hDDDD	;
				14'b11110101000001: Data_out <= 16'hDDE9	;
				14'b11110101000010: Data_out <= 16'hDDF5	;
				14'b11110101000011: Data_out <= 16'hDE01	;
				14'b11110101000100: Data_out <= 16'hDE0D	;
				14'b11110101000101: Data_out <= 16'hDE19	;
				14'b11110101000110: Data_out <= 16'hDE25	;
				14'b11110101000111: Data_out <= 16'hDE32	;
				14'b11110101001000: Data_out <= 16'hDE3E	;
				14'b11110101001001: Data_out <= 16'hDE4A	;
				14'b11110101001010: Data_out <= 16'hDE56	;
				14'b11110101001011: Data_out <= 16'hDE62	;
				14'b11110101001100: Data_out <= 16'hDE6E	;
				14'b11110101001101: Data_out <= 16'hDE7A	;
				14'b11110101001110: Data_out <= 16'hDE86	;
				14'b11110101001111: Data_out <= 16'hDE93	;
				14'b11110101010000: Data_out <= 16'hDE9F	;
				14'b11110101010001: Data_out <= 16'hDEAB	;
				14'b11110101010010: Data_out <= 16'hDEB7	;
				14'b11110101010011: Data_out <= 16'hDEC3	;
				14'b11110101010100: Data_out <= 16'hDECF	;
				14'b11110101010101: Data_out <= 16'hDEDB	;
				14'b11110101010110: Data_out <= 16'hDEE7	;
				14'b11110101010111: Data_out <= 16'hDEF4	;
				14'b11110101011000: Data_out <= 16'hDF00	;
				14'b11110101011001: Data_out <= 16'hDF0C	;
				14'b11110101011010: Data_out <= 16'hDF18	;
				14'b11110101011011: Data_out <= 16'hDF24	;
				14'b11110101011100: Data_out <= 16'hDF30	;
				14'b11110101011101: Data_out <= 16'hDF3C	;
				14'b11110101011110: Data_out <= 16'hDF49	;
				14'b11110101011111: Data_out <= 16'hDF55	;
				14'b11110101100000: Data_out <= 16'hDF61	;
				14'b11110101100001: Data_out <= 16'hDF6D	;
				14'b11110101100010: Data_out <= 16'hDF79	;
				14'b11110101100011: Data_out <= 16'hDF85	;
				14'b11110101100100: Data_out <= 16'hDF92	;
				14'b11110101100101: Data_out <= 16'hDF9E	;
				14'b11110101100110: Data_out <= 16'hDFAA	;
				14'b11110101100111: Data_out <= 16'hDFB6	;
				14'b11110101101000: Data_out <= 16'hDFC2	;
				14'b11110101101001: Data_out <= 16'hDFCE	;
				14'b11110101101010: Data_out <= 16'hDFDA	;
				14'b11110101101011: Data_out <= 16'hDFE7	;
				14'b11110101101100: Data_out <= 16'hDFF3	;
				14'b11110101101101: Data_out <= 16'hDFFF	;
				14'b11110101101110: Data_out <= 16'hE00B	;
				14'b11110101101111: Data_out <= 16'hE017	;
				14'b11110101110000: Data_out <= 16'hE023	;
				14'b11110101110001: Data_out <= 16'hE030	;
				14'b11110101110010: Data_out <= 16'hE03C	;
				14'b11110101110011: Data_out <= 16'hE048	;
				14'b11110101110100: Data_out <= 16'hE054	;
				14'b11110101110101: Data_out <= 16'hE060	;
				14'b11110101110110: Data_out <= 16'hE06D	;
				14'b11110101110111: Data_out <= 16'hE079	;
				14'b11110101111000: Data_out <= 16'hE085	;
				14'b11110101111001: Data_out <= 16'hE091	;
				14'b11110101111010: Data_out <= 16'hE09D	;
				14'b11110101111011: Data_out <= 16'hE0A9	;
				14'b11110101111100: Data_out <= 16'hE0B6	;
				14'b11110101111101: Data_out <= 16'hE0C2	;
				14'b11110101111110: Data_out <= 16'hE0CE	;
				14'b11110101111111: Data_out <= 16'hE0DA	;
				14'b11110110000000: Data_out <= 16'hE0E6	;
				14'b11110110000001: Data_out <= 16'hE0F3	;
				14'b11110110000010: Data_out <= 16'hE0FF	;
				14'b11110110000011: Data_out <= 16'hE10B	;
				14'b11110110000100: Data_out <= 16'hE117	;
				14'b11110110000101: Data_out <= 16'hE123	;
				14'b11110110000110: Data_out <= 16'hE130	;
				14'b11110110000111: Data_out <= 16'hE13C	;
				14'b11110110001000: Data_out <= 16'hE148	;
				14'b11110110001001: Data_out <= 16'hE154	;
				14'b11110110001010: Data_out <= 16'hE160	;
				14'b11110110001011: Data_out <= 16'hE16D	;
				14'b11110110001100: Data_out <= 16'hE179	;
				14'b11110110001101: Data_out <= 16'hE185	;
				14'b11110110001110: Data_out <= 16'hE191	;
				14'b11110110001111: Data_out <= 16'hE19D	;
				14'b11110110010000: Data_out <= 16'hE1AA	;
				14'b11110110010001: Data_out <= 16'hE1B6	;
				14'b11110110010010: Data_out <= 16'hE1C2	;
				14'b11110110010011: Data_out <= 16'hE1CE	;
				14'b11110110010100: Data_out <= 16'hE1DA	;
				14'b11110110010101: Data_out <= 16'hE1E7	;
				14'b11110110010110: Data_out <= 16'hE1F3	;
				14'b11110110010111: Data_out <= 16'hE1FF	;
				14'b11110110011000: Data_out <= 16'hE20B	;
				14'b11110110011001: Data_out <= 16'hE217	;
				14'b11110110011010: Data_out <= 16'hE224	;
				14'b11110110011011: Data_out <= 16'hE230	;
				14'b11110110011100: Data_out <= 16'hE23C	;
				14'b11110110011101: Data_out <= 16'hE248	;
				14'b11110110011110: Data_out <= 16'hE255	;
				14'b11110110011111: Data_out <= 16'hE261	;
				14'b11110110100000: Data_out <= 16'hE26D	;
				14'b11110110100001: Data_out <= 16'hE279	;
				14'b11110110100010: Data_out <= 16'hE285	;
				14'b11110110100011: Data_out <= 16'hE292	;
				14'b11110110100100: Data_out <= 16'hE29E	;
				14'b11110110100101: Data_out <= 16'hE2AA	;
				14'b11110110100110: Data_out <= 16'hE2B6	;
				14'b11110110100111: Data_out <= 16'hE2C3	;
				14'b11110110101000: Data_out <= 16'hE2CF	;
				14'b11110110101001: Data_out <= 16'hE2DB	;
				14'b11110110101010: Data_out <= 16'hE2E7	;
				14'b11110110101011: Data_out <= 16'hE2F4	;
				14'b11110110101100: Data_out <= 16'hE300	;
				14'b11110110101101: Data_out <= 16'hE30C	;
				14'b11110110101110: Data_out <= 16'hE318	;
				14'b11110110101111: Data_out <= 16'hE325	;
				14'b11110110110000: Data_out <= 16'hE331	;
				14'b11110110110001: Data_out <= 16'hE33D	;
				14'b11110110110010: Data_out <= 16'hE349	;
				14'b11110110110011: Data_out <= 16'hE356	;
				14'b11110110110100: Data_out <= 16'hE362	;
				14'b11110110110101: Data_out <= 16'hE36E	;
				14'b11110110110110: Data_out <= 16'hE37A	;
				14'b11110110110111: Data_out <= 16'hE387	;
				14'b11110110111000: Data_out <= 16'hE393	;
				14'b11110110111001: Data_out <= 16'hE39F	;
				14'b11110110111010: Data_out <= 16'hE3AB	;
				14'b11110110111011: Data_out <= 16'hE3B8	;
				14'b11110110111100: Data_out <= 16'hE3C4	;
				14'b11110110111101: Data_out <= 16'hE3D0	;
				14'b11110110111110: Data_out <= 16'hE3DC	;
				14'b11110110111111: Data_out <= 16'hE3E9	;
				14'b11110111000000: Data_out <= 16'hE3F5	;
				14'b11110111000001: Data_out <= 16'hE401	;
				14'b11110111000010: Data_out <= 16'hE40D	;
				14'b11110111000011: Data_out <= 16'hE41A	;
				14'b11110111000100: Data_out <= 16'hE426	;
				14'b11110111000101: Data_out <= 16'hE432	;
				14'b11110111000110: Data_out <= 16'hE43E	;
				14'b11110111000111: Data_out <= 16'hE44B	;
				14'b11110111001000: Data_out <= 16'hE457	;
				14'b11110111001001: Data_out <= 16'hE463	;
				14'b11110111001010: Data_out <= 16'hE46F	;
				14'b11110111001011: Data_out <= 16'hE47C	;
				14'b11110111001100: Data_out <= 16'hE488	;
				14'b11110111001101: Data_out <= 16'hE494	;
				14'b11110111001110: Data_out <= 16'hE4A1	;
				14'b11110111001111: Data_out <= 16'hE4AD	;
				14'b11110111010000: Data_out <= 16'hE4B9	;
				14'b11110111010001: Data_out <= 16'hE4C5	;
				14'b11110111010010: Data_out <= 16'hE4D2	;
				14'b11110111010011: Data_out <= 16'hE4DE	;
				14'b11110111010100: Data_out <= 16'hE4EA	;
				14'b11110111010101: Data_out <= 16'hE4F7	;
				14'b11110111010110: Data_out <= 16'hE503	;
				14'b11110111010111: Data_out <= 16'hE50F	;
				14'b11110111011000: Data_out <= 16'hE51B	;
				14'b11110111011001: Data_out <= 16'hE528	;
				14'b11110111011010: Data_out <= 16'hE534	;
				14'b11110111011011: Data_out <= 16'hE540	;
				14'b11110111011100: Data_out <= 16'hE54D	;
				14'b11110111011101: Data_out <= 16'hE559	;
				14'b11110111011110: Data_out <= 16'hE565	;
				14'b11110111011111: Data_out <= 16'hE571	;
				14'b11110111100000: Data_out <= 16'hE57E	;
				14'b11110111100001: Data_out <= 16'hE58A	;
				14'b11110111100010: Data_out <= 16'hE596	;
				14'b11110111100011: Data_out <= 16'hE5A3	;
				14'b11110111100100: Data_out <= 16'hE5AF	;
				14'b11110111100101: Data_out <= 16'hE5BB	;
				14'b11110111100110: Data_out <= 16'hE5C7	;
				14'b11110111100111: Data_out <= 16'hE5D4	;
				14'b11110111101000: Data_out <= 16'hE5E0	;
				14'b11110111101001: Data_out <= 16'hE5EC	;
				14'b11110111101010: Data_out <= 16'hE5F9	;
				14'b11110111101011: Data_out <= 16'hE605	;
				14'b11110111101100: Data_out <= 16'hE611	;
				14'b11110111101101: Data_out <= 16'hE61E	;
				14'b11110111101110: Data_out <= 16'hE62A	;
				14'b11110111101111: Data_out <= 16'hE636	;
				14'b11110111110000: Data_out <= 16'hE643	;
				14'b11110111110001: Data_out <= 16'hE64F	;
				14'b11110111110010: Data_out <= 16'hE65B	;
				14'b11110111110011: Data_out <= 16'hE667	;
				14'b11110111110100: Data_out <= 16'hE674	;
				14'b11110111110101: Data_out <= 16'hE680	;
				14'b11110111110110: Data_out <= 16'hE68C	;
				14'b11110111110111: Data_out <= 16'hE699	;
				14'b11110111111000: Data_out <= 16'hE6A5	;
				14'b11110111111001: Data_out <= 16'hE6B1	;
				14'b11110111111010: Data_out <= 16'hE6BE	;
				14'b11110111111011: Data_out <= 16'hE6CA	;
				14'b11110111111100: Data_out <= 16'hE6D6	;
				14'b11110111111101: Data_out <= 16'hE6E3	;
				14'b11110111111110: Data_out <= 16'hE6EF	;
				14'b11110111111111: Data_out <= 16'hE6FB	;
				14'b11111000000000: Data_out <= 16'hE708	;
				14'b11111000000001: Data_out <= 16'hE714	;
				14'b11111000000010: Data_out <= 16'hE720	;
				14'b11111000000011: Data_out <= 16'hE72D	;
				14'b11111000000100: Data_out <= 16'hE739	;
				14'b11111000000101: Data_out <= 16'hE745	;
				14'b11111000000110: Data_out <= 16'hE752	;
				14'b11111000000111: Data_out <= 16'hE75E	;
				14'b11111000001000: Data_out <= 16'hE76A	;
				14'b11111000001001: Data_out <= 16'hE777	;
				14'b11111000001010: Data_out <= 16'hE783	;
				14'b11111000001011: Data_out <= 16'hE78F	;
				14'b11111000001100: Data_out <= 16'hE79C	;
				14'b11111000001101: Data_out <= 16'hE7A8	;
				14'b11111000001110: Data_out <= 16'hE7B4	;
				14'b11111000001111: Data_out <= 16'hE7C1	;
				14'b11111000010000: Data_out <= 16'hE7CD	;
				14'b11111000010001: Data_out <= 16'hE7D9	;
				14'b11111000010010: Data_out <= 16'hE7E6	;
				14'b11111000010011: Data_out <= 16'hE7F2	;
				14'b11111000010100: Data_out <= 16'hE7FE	;
				14'b11111000010101: Data_out <= 16'hE80B	;
				14'b11111000010110: Data_out <= 16'hE817	;
				14'b11111000010111: Data_out <= 16'hE823	;
				14'b11111000011000: Data_out <= 16'hE830	;
				14'b11111000011001: Data_out <= 16'hE83C	;
				14'b11111000011010: Data_out <= 16'hE848	;
				14'b11111000011011: Data_out <= 16'hE855	;
				14'b11111000011100: Data_out <= 16'hE861	;
				14'b11111000011101: Data_out <= 16'hE86D	;
				14'b11111000011110: Data_out <= 16'hE87A	;
				14'b11111000011111: Data_out <= 16'hE886	;
				14'b11111000100000: Data_out <= 16'hE892	;
				14'b11111000100001: Data_out <= 16'hE89F	;
				14'b11111000100010: Data_out <= 16'hE8AB	;
				14'b11111000100011: Data_out <= 16'hE8B7	;
				14'b11111000100100: Data_out <= 16'hE8C4	;
				14'b11111000100101: Data_out <= 16'hE8D0	;
				14'b11111000100110: Data_out <= 16'hE8DD	;
				14'b11111000100111: Data_out <= 16'hE8E9	;
				14'b11111000101000: Data_out <= 16'hE8F5	;
				14'b11111000101001: Data_out <= 16'hE902	;
				14'b11111000101010: Data_out <= 16'hE90E	;
				14'b11111000101011: Data_out <= 16'hE91A	;
				14'b11111000101100: Data_out <= 16'hE927	;
				14'b11111000101101: Data_out <= 16'hE933	;
				14'b11111000101110: Data_out <= 16'hE93F	;
				14'b11111000101111: Data_out <= 16'hE94C	;
				14'b11111000110000: Data_out <= 16'hE958	;
				14'b11111000110001: Data_out <= 16'hE965	;
				14'b11111000110010: Data_out <= 16'hE971	;
				14'b11111000110011: Data_out <= 16'hE97D	;
				14'b11111000110100: Data_out <= 16'hE98A	;
				14'b11111000110101: Data_out <= 16'hE996	;
				14'b11111000110110: Data_out <= 16'hE9A2	;
				14'b11111000110111: Data_out <= 16'hE9AF	;
				14'b11111000111000: Data_out <= 16'hE9BB	;
				14'b11111000111001: Data_out <= 16'hE9C8	;
				14'b11111000111010: Data_out <= 16'hE9D4	;
				14'b11111000111011: Data_out <= 16'hE9E0	;
				14'b11111000111100: Data_out <= 16'hE9ED	;
				14'b11111000111101: Data_out <= 16'hE9F9	;
				14'b11111000111110: Data_out <= 16'hEA05	;
				14'b11111000111111: Data_out <= 16'hEA12	;
				14'b11111001000000: Data_out <= 16'hEA1E	;
				14'b11111001000001: Data_out <= 16'hEA2B	;
				14'b11111001000010: Data_out <= 16'hEA37	;
				14'b11111001000011: Data_out <= 16'hEA43	;
				14'b11111001000100: Data_out <= 16'hEA50	;
				14'b11111001000101: Data_out <= 16'hEA5C	;
				14'b11111001000110: Data_out <= 16'hEA68	;
				14'b11111001000111: Data_out <= 16'hEA75	;
				14'b11111001001000: Data_out <= 16'hEA81	;
				14'b11111001001001: Data_out <= 16'hEA8E	;
				14'b11111001001010: Data_out <= 16'hEA9A	;
				14'b11111001001011: Data_out <= 16'hEAA6	;
				14'b11111001001100: Data_out <= 16'hEAB3	;
				14'b11111001001101: Data_out <= 16'hEABF	;
				14'b11111001001110: Data_out <= 16'hEACC	;
				14'b11111001001111: Data_out <= 16'hEAD8	;
				14'b11111001010000: Data_out <= 16'hEAE4	;
				14'b11111001010001: Data_out <= 16'hEAF1	;
				14'b11111001010010: Data_out <= 16'hEAFD	;
				14'b11111001010011: Data_out <= 16'hEB0A	;
				14'b11111001010100: Data_out <= 16'hEB16	;
				14'b11111001010101: Data_out <= 16'hEB22	;
				14'b11111001010110: Data_out <= 16'hEB2F	;
				14'b11111001010111: Data_out <= 16'hEB3B	;
				14'b11111001011000: Data_out <= 16'hEB48	;
				14'b11111001011001: Data_out <= 16'hEB54	;
				14'b11111001011010: Data_out <= 16'hEB60	;
				14'b11111001011011: Data_out <= 16'hEB6D	;
				14'b11111001011100: Data_out <= 16'hEB79	;
				14'b11111001011101: Data_out <= 16'hEB86	;
				14'b11111001011110: Data_out <= 16'hEB92	;
				14'b11111001011111: Data_out <= 16'hEB9E	;
				14'b11111001100000: Data_out <= 16'hEBAB	;
				14'b11111001100001: Data_out <= 16'hEBB7	;
				14'b11111001100010: Data_out <= 16'hEBC4	;
				14'b11111001100011: Data_out <= 16'hEBD0	;
				14'b11111001100100: Data_out <= 16'hEBDC	;
				14'b11111001100101: Data_out <= 16'hEBE9	;
				14'b11111001100110: Data_out <= 16'hEBF5	;
				14'b11111001100111: Data_out <= 16'hEC02	;
				14'b11111001101000: Data_out <= 16'hEC0E	;
				14'b11111001101001: Data_out <= 16'hEC1A	;
				14'b11111001101010: Data_out <= 16'hEC27	;
				14'b11111001101011: Data_out <= 16'hEC33	;
				14'b11111001101100: Data_out <= 16'hEC40	;
				14'b11111001101101: Data_out <= 16'hEC4C	;
				14'b11111001101110: Data_out <= 16'hEC59	;
				14'b11111001101111: Data_out <= 16'hEC65	;
				14'b11111001110000: Data_out <= 16'hEC71	;
				14'b11111001110001: Data_out <= 16'hEC7E	;
				14'b11111001110010: Data_out <= 16'hEC8A	;
				14'b11111001110011: Data_out <= 16'hEC97	;
				14'b11111001110100: Data_out <= 16'hECA3	;
				14'b11111001110101: Data_out <= 16'hECAF	;
				14'b11111001110110: Data_out <= 16'hECBC	;
				14'b11111001110111: Data_out <= 16'hECC8	;
				14'b11111001111000: Data_out <= 16'hECD5	;
				14'b11111001111001: Data_out <= 16'hECE1	;
				14'b11111001111010: Data_out <= 16'hECEE	;
				14'b11111001111011: Data_out <= 16'hECFA	;
				14'b11111001111100: Data_out <= 16'hED06	;
				14'b11111001111101: Data_out <= 16'hED13	;
				14'b11111001111110: Data_out <= 16'hED1F	;
				14'b11111001111111: Data_out <= 16'hED2C	;
				14'b11111010000000: Data_out <= 16'hED38	;
				14'b11111010000001: Data_out <= 16'hED45	;
				14'b11111010000010: Data_out <= 16'hED51	;
				14'b11111010000011: Data_out <= 16'hED5D	;
				14'b11111010000100: Data_out <= 16'hED6A	;
				14'b11111010000101: Data_out <= 16'hED76	;
				14'b11111010000110: Data_out <= 16'hED83	;
				14'b11111010000111: Data_out <= 16'hED8F	;
				14'b11111010001000: Data_out <= 16'hED9C	;
				14'b11111010001001: Data_out <= 16'hEDA8	;
				14'b11111010001010: Data_out <= 16'hEDB5	;
				14'b11111010001011: Data_out <= 16'hEDC1	;
				14'b11111010001100: Data_out <= 16'hEDCD	;
				14'b11111010001101: Data_out <= 16'hEDDA	;
				14'b11111010001110: Data_out <= 16'hEDE6	;
				14'b11111010001111: Data_out <= 16'hEDF3	;
				14'b11111010010000: Data_out <= 16'hEDFF	;
				14'b11111010010001: Data_out <= 16'hEE0C	;
				14'b11111010010010: Data_out <= 16'hEE18	;
				14'b11111010010011: Data_out <= 16'hEE24	;
				14'b11111010010100: Data_out <= 16'hEE31	;
				14'b11111010010101: Data_out <= 16'hEE3D	;
				14'b11111010010110: Data_out <= 16'hEE4A	;
				14'b11111010010111: Data_out <= 16'hEE56	;
				14'b11111010011000: Data_out <= 16'hEE63	;
				14'b11111010011001: Data_out <= 16'hEE6F	;
				14'b11111010011010: Data_out <= 16'hEE7C	;
				14'b11111010011011: Data_out <= 16'hEE88	;
				14'b11111010011100: Data_out <= 16'hEE94	;
				14'b11111010011101: Data_out <= 16'hEEA1	;
				14'b11111010011110: Data_out <= 16'hEEAD	;
				14'b11111010011111: Data_out <= 16'hEEBA	;
				14'b11111010100000: Data_out <= 16'hEEC6	;
				14'b11111010100001: Data_out <= 16'hEED3	;
				14'b11111010100010: Data_out <= 16'hEEDF	;
				14'b11111010100011: Data_out <= 16'hEEEC	;
				14'b11111010100100: Data_out <= 16'hEEF8	;
				14'b11111010100101: Data_out <= 16'hEF05	;
				14'b11111010100110: Data_out <= 16'hEF11	;
				14'b11111010100111: Data_out <= 16'hEF1D	;
				14'b11111010101000: Data_out <= 16'hEF2A	;
				14'b11111010101001: Data_out <= 16'hEF36	;
				14'b11111010101010: Data_out <= 16'hEF43	;
				14'b11111010101011: Data_out <= 16'hEF4F	;
				14'b11111010101100: Data_out <= 16'hEF5C	;
				14'b11111010101101: Data_out <= 16'hEF68	;
				14'b11111010101110: Data_out <= 16'hEF75	;
				14'b11111010101111: Data_out <= 16'hEF81	;
				14'b11111010110000: Data_out <= 16'hEF8E	;
				14'b11111010110001: Data_out <= 16'hEF9A	;
				14'b11111010110010: Data_out <= 16'hEFA7	;
				14'b11111010110011: Data_out <= 16'hEFB3	;
				14'b11111010110100: Data_out <= 16'hEFBF	;
				14'b11111010110101: Data_out <= 16'hEFCC	;
				14'b11111010110110: Data_out <= 16'hEFD8	;
				14'b11111010110111: Data_out <= 16'hEFE5	;
				14'b11111010111000: Data_out <= 16'hEFF1	;
				14'b11111010111001: Data_out <= 16'hEFFE	;
				14'b11111010111010: Data_out <= 16'hF00A	;
				14'b11111010111011: Data_out <= 16'hF017	;
				14'b11111010111100: Data_out <= 16'hF023	;
				14'b11111010111101: Data_out <= 16'hF030	;
				14'b11111010111110: Data_out <= 16'hF03C	;
				14'b11111010111111: Data_out <= 16'hF049	;
				14'b11111011000000: Data_out <= 16'hF055	;
				14'b11111011000001: Data_out <= 16'hF062	;
				14'b11111011000010: Data_out <= 16'hF06E	;
				14'b11111011000011: Data_out <= 16'hF07A	;
				14'b11111011000100: Data_out <= 16'hF087	;
				14'b11111011000101: Data_out <= 16'hF093	;
				14'b11111011000110: Data_out <= 16'hF0A0	;
				14'b11111011000111: Data_out <= 16'hF0AC	;
				14'b11111011001000: Data_out <= 16'hF0B9	;
				14'b11111011001001: Data_out <= 16'hF0C5	;
				14'b11111011001010: Data_out <= 16'hF0D2	;
				14'b11111011001011: Data_out <= 16'hF0DE	;
				14'b11111011001100: Data_out <= 16'hF0EB	;
				14'b11111011001101: Data_out <= 16'hF0F7	;
				14'b11111011001110: Data_out <= 16'hF104	;
				14'b11111011001111: Data_out <= 16'hF110	;
				14'b11111011010000: Data_out <= 16'hF11D	;
				14'b11111011010001: Data_out <= 16'hF129	;
				14'b11111011010010: Data_out <= 16'hF136	;
				14'b11111011010011: Data_out <= 16'hF142	;
				14'b11111011010100: Data_out <= 16'hF14F	;
				14'b11111011010101: Data_out <= 16'hF15B	;
				14'b11111011010110: Data_out <= 16'hF168	;
				14'b11111011010111: Data_out <= 16'hF174	;
				14'b11111011011000: Data_out <= 16'hF181	;
				14'b11111011011001: Data_out <= 16'hF18D	;
				14'b11111011011010: Data_out <= 16'hF19A	;
				14'b11111011011011: Data_out <= 16'hF1A6	;
				14'b11111011011100: Data_out <= 16'hF1B2	;
				14'b11111011011101: Data_out <= 16'hF1BF	;
				14'b11111011011110: Data_out <= 16'hF1CB	;
				14'b11111011011111: Data_out <= 16'hF1D8	;
				14'b11111011100000: Data_out <= 16'hF1E4	;
				14'b11111011100001: Data_out <= 16'hF1F1	;
				14'b11111011100010: Data_out <= 16'hF1FD	;
				14'b11111011100011: Data_out <= 16'hF20A	;
				14'b11111011100100: Data_out <= 16'hF216	;
				14'b11111011100101: Data_out <= 16'hF223	;
				14'b11111011100110: Data_out <= 16'hF22F	;
				14'b11111011100111: Data_out <= 16'hF23C	;
				14'b11111011101000: Data_out <= 16'hF248	;
				14'b11111011101001: Data_out <= 16'hF255	;
				14'b11111011101010: Data_out <= 16'hF261	;
				14'b11111011101011: Data_out <= 16'hF26E	;
				14'b11111011101100: Data_out <= 16'hF27A	;
				14'b11111011101101: Data_out <= 16'hF287	;
				14'b11111011101110: Data_out <= 16'hF293	;
				14'b11111011101111: Data_out <= 16'hF2A0	;
				14'b11111011110000: Data_out <= 16'hF2AC	;
				14'b11111011110001: Data_out <= 16'hF2B9	;
				14'b11111011110010: Data_out <= 16'hF2C5	;
				14'b11111011110011: Data_out <= 16'hF2D2	;
				14'b11111011110100: Data_out <= 16'hF2DE	;
				14'b11111011110101: Data_out <= 16'hF2EB	;
				14'b11111011110110: Data_out <= 16'hF2F7	;
				14'b11111011110111: Data_out <= 16'hF304	;
				14'b11111011111000: Data_out <= 16'hF310	;
				14'b11111011111001: Data_out <= 16'hF31D	;
				14'b11111011111010: Data_out <= 16'hF329	;
				14'b11111011111011: Data_out <= 16'hF336	;
				14'b11111011111100: Data_out <= 16'hF342	;
				14'b11111011111101: Data_out <= 16'hF34F	;
				14'b11111011111110: Data_out <= 16'hF35B	;
				14'b11111011111111: Data_out <= 16'hF368	;
				14'b11111100000000: Data_out <= 16'hF374	;
				14'b11111100000001: Data_out <= 16'hF381	;
				14'b11111100000010: Data_out <= 16'hF38D	;
				14'b11111100000011: Data_out <= 16'hF39A	;
				14'b11111100000100: Data_out <= 16'hF3A6	;
				14'b11111100000101: Data_out <= 16'hF3B3	;
				14'b11111100000110: Data_out <= 16'hF3BF	;
				14'b11111100000111: Data_out <= 16'hF3CC	;
				14'b11111100001000: Data_out <= 16'hF3D8	;
				14'b11111100001001: Data_out <= 16'hF3E5	;
				14'b11111100001010: Data_out <= 16'hF3F1	;
				14'b11111100001011: Data_out <= 16'hF3FE	;
				14'b11111100001100: Data_out <= 16'hF40A	;
				14'b11111100001101: Data_out <= 16'hF417	;
				14'b11111100001110: Data_out <= 16'hF423	;
				14'b11111100001111: Data_out <= 16'hF430	;
				14'b11111100010000: Data_out <= 16'hF43D	;
				14'b11111100010001: Data_out <= 16'hF449	;
				14'b11111100010010: Data_out <= 16'hF456	;
				14'b11111100010011: Data_out <= 16'hF462	;
				14'b11111100010100: Data_out <= 16'hF46F	;
				14'b11111100010101: Data_out <= 16'hF47B	;
				14'b11111100010110: Data_out <= 16'hF488	;
				14'b11111100010111: Data_out <= 16'hF494	;
				14'b11111100011000: Data_out <= 16'hF4A1	;
				14'b11111100011001: Data_out <= 16'hF4AD	;
				14'b11111100011010: Data_out <= 16'hF4BA	;
				14'b11111100011011: Data_out <= 16'hF4C6	;
				14'b11111100011100: Data_out <= 16'hF4D3	;
				14'b11111100011101: Data_out <= 16'hF4DF	;
				14'b11111100011110: Data_out <= 16'hF4EC	;
				14'b11111100011111: Data_out <= 16'hF4F8	;
				14'b11111100100000: Data_out <= 16'hF505	;
				14'b11111100100001: Data_out <= 16'hF511	;
				14'b11111100100010: Data_out <= 16'hF51E	;
				14'b11111100100011: Data_out <= 16'hF52A	;
				14'b11111100100100: Data_out <= 16'hF537	;
				14'b11111100100101: Data_out <= 16'hF543	;
				14'b11111100100110: Data_out <= 16'hF550	;
				14'b11111100100111: Data_out <= 16'hF55C	;
				14'b11111100101000: Data_out <= 16'hF569	;
				14'b11111100101001: Data_out <= 16'hF575	;
				14'b11111100101010: Data_out <= 16'hF582	;
				14'b11111100101011: Data_out <= 16'hF58F	;
				14'b11111100101100: Data_out <= 16'hF59B	;
				14'b11111100101101: Data_out <= 16'hF5A8	;
				14'b11111100101110: Data_out <= 16'hF5B4	;
				14'b11111100101111: Data_out <= 16'hF5C1	;
				14'b11111100110000: Data_out <= 16'hF5CD	;
				14'b11111100110001: Data_out <= 16'hF5DA	;
				14'b11111100110010: Data_out <= 16'hF5E6	;
				14'b11111100110011: Data_out <= 16'hF5F3	;
				14'b11111100110100: Data_out <= 16'hF5FF	;
				14'b11111100110101: Data_out <= 16'hF60C	;
				14'b11111100110110: Data_out <= 16'hF618	;
				14'b11111100110111: Data_out <= 16'hF625	;
				14'b11111100111000: Data_out <= 16'hF631	;
				14'b11111100111001: Data_out <= 16'hF63E	;
				14'b11111100111010: Data_out <= 16'hF64A	;
				14'b11111100111011: Data_out <= 16'hF657	;
				14'b11111100111100: Data_out <= 16'hF663	;
				14'b11111100111101: Data_out <= 16'hF670	;
				14'b11111100111110: Data_out <= 16'hF67D	;
				14'b11111100111111: Data_out <= 16'hF689	;
				14'b11111101000000: Data_out <= 16'hF696	;
				14'b11111101000001: Data_out <= 16'hF6A2	;
				14'b11111101000010: Data_out <= 16'hF6AF	;
				14'b11111101000011: Data_out <= 16'hF6BB	;
				14'b11111101000100: Data_out <= 16'hF6C8	;
				14'b11111101000101: Data_out <= 16'hF6D4	;
				14'b11111101000110: Data_out <= 16'hF6E1	;
				14'b11111101000111: Data_out <= 16'hF6ED	;
				14'b11111101001000: Data_out <= 16'hF6FA	;
				14'b11111101001001: Data_out <= 16'hF706	;
				14'b11111101001010: Data_out <= 16'hF713	;
				14'b11111101001011: Data_out <= 16'hF71F	;
				14'b11111101001100: Data_out <= 16'hF72C	;
				14'b11111101001101: Data_out <= 16'hF739	;
				14'b11111101001110: Data_out <= 16'hF745	;
				14'b11111101001111: Data_out <= 16'hF752	;
				14'b11111101010000: Data_out <= 16'hF75E	;
				14'b11111101010001: Data_out <= 16'hF76B	;
				14'b11111101010010: Data_out <= 16'hF777	;
				14'b11111101010011: Data_out <= 16'hF784	;
				14'b11111101010100: Data_out <= 16'hF790	;
				14'b11111101010101: Data_out <= 16'hF79D	;
				14'b11111101010110: Data_out <= 16'hF7A9	;
				14'b11111101010111: Data_out <= 16'hF7B6	;
				14'b11111101011000: Data_out <= 16'hF7C2	;
				14'b11111101011001: Data_out <= 16'hF7CF	;
				14'b11111101011010: Data_out <= 16'hF7DC	;
				14'b11111101011011: Data_out <= 16'hF7E8	;
				14'b11111101011100: Data_out <= 16'hF7F5	;
				14'b11111101011101: Data_out <= 16'hF801	;
				14'b11111101011110: Data_out <= 16'hF80E	;
				14'b11111101011111: Data_out <= 16'hF81A	;
				14'b11111101100000: Data_out <= 16'hF827	;
				14'b11111101100001: Data_out <= 16'hF833	;
				14'b11111101100010: Data_out <= 16'hF840	;
				14'b11111101100011: Data_out <= 16'hF84C	;
				14'b11111101100100: Data_out <= 16'hF859	;
				14'b11111101100101: Data_out <= 16'hF866	;
				14'b11111101100110: Data_out <= 16'hF872	;
				14'b11111101100111: Data_out <= 16'hF87F	;
				14'b11111101101000: Data_out <= 16'hF88B	;
				14'b11111101101001: Data_out <= 16'hF898	;
				14'b11111101101010: Data_out <= 16'hF8A4	;
				14'b11111101101011: Data_out <= 16'hF8B1	;
				14'b11111101101100: Data_out <= 16'hF8BD	;
				14'b11111101101101: Data_out <= 16'hF8CA	;
				14'b11111101101110: Data_out <= 16'hF8D6	;
				14'b11111101101111: Data_out <= 16'hF8E3	;
				14'b11111101110000: Data_out <= 16'hF8F0	;
				14'b11111101110001: Data_out <= 16'hF8FC	;
				14'b11111101110010: Data_out <= 16'hF909	;
				14'b11111101110011: Data_out <= 16'hF915	;
				14'b11111101110100: Data_out <= 16'hF922	;
				14'b11111101110101: Data_out <= 16'hF92E	;
				14'b11111101110110: Data_out <= 16'hF93B	;
				14'b11111101110111: Data_out <= 16'hF947	;
				14'b11111101111000: Data_out <= 16'hF954	;
				14'b11111101111001: Data_out <= 16'hF960	;
				14'b11111101111010: Data_out <= 16'hF96D	;
				14'b11111101111011: Data_out <= 16'hF97A	;
				14'b11111101111100: Data_out <= 16'hF986	;
				14'b11111101111101: Data_out <= 16'hF993	;
				14'b11111101111110: Data_out <= 16'hF99F	;
				14'b11111101111111: Data_out <= 16'hF9AC	;
				14'b11111110000000: Data_out <= 16'hF9B8	;
				14'b11111110000001: Data_out <= 16'hF9C5	;
				14'b11111110000010: Data_out <= 16'hF9D1	;
				14'b11111110000011: Data_out <= 16'hF9DE	;
				14'b11111110000100: Data_out <= 16'hF9EB	;
				14'b11111110000101: Data_out <= 16'hF9F7	;
				14'b11111110000110: Data_out <= 16'hFA04	;
				14'b11111110000111: Data_out <= 16'hFA10	;
				14'b11111110001000: Data_out <= 16'hFA1D	;
				14'b11111110001001: Data_out <= 16'hFA29	;
				14'b11111110001010: Data_out <= 16'hFA36	;
				14'b11111110001011: Data_out <= 16'hFA42	;
				14'b11111110001100: Data_out <= 16'hFA4F	;
				14'b11111110001101: Data_out <= 16'hFA5B	;
				14'b11111110001110: Data_out <= 16'hFA68	;
				14'b11111110001111: Data_out <= 16'hFA75	;
				14'b11111110010000: Data_out <= 16'hFA81	;
				14'b11111110010001: Data_out <= 16'hFA8E	;
				14'b11111110010010: Data_out <= 16'hFA9A	;
				14'b11111110010011: Data_out <= 16'hFAA7	;
				14'b11111110010100: Data_out <= 16'hFAB3	;
				14'b11111110010101: Data_out <= 16'hFAC0	;
				14'b11111110010110: Data_out <= 16'hFACC	;
				14'b11111110010111: Data_out <= 16'hFAD9	;
				14'b11111110011000: Data_out <= 16'hFAE6	;
				14'b11111110011001: Data_out <= 16'hFAF2	;
				14'b11111110011010: Data_out <= 16'hFAFF	;
				14'b11111110011011: Data_out <= 16'hFB0B	;
				14'b11111110011100: Data_out <= 16'hFB18	;
				14'b11111110011101: Data_out <= 16'hFB24	;
				14'b11111110011110: Data_out <= 16'hFB31	;
				14'b11111110011111: Data_out <= 16'hFB3D	;
				14'b11111110100000: Data_out <= 16'hFB4A	;
				14'b11111110100001: Data_out <= 16'hFB57	;
				14'b11111110100010: Data_out <= 16'hFB63	;
				14'b11111110100011: Data_out <= 16'hFB70	;
				14'b11111110100100: Data_out <= 16'hFB7C	;
				14'b11111110100101: Data_out <= 16'hFB89	;
				14'b11111110100110: Data_out <= 16'hFB95	;
				14'b11111110100111: Data_out <= 16'hFBA2	;
				14'b11111110101000: Data_out <= 16'hFBAF	;
				14'b11111110101001: Data_out <= 16'hFBBB	;
				14'b11111110101010: Data_out <= 16'hFBC8	;
				14'b11111110101011: Data_out <= 16'hFBD4	;
				14'b11111110101100: Data_out <= 16'hFBE1	;
				14'b11111110101101: Data_out <= 16'hFBED	;
				14'b11111110101110: Data_out <= 16'hFBFA	;
				14'b11111110101111: Data_out <= 16'hFC06	;
				14'b11111110110000: Data_out <= 16'hFC13	;
				14'b11111110110001: Data_out <= 16'hFC20	;
				14'b11111110110010: Data_out <= 16'hFC2C	;
				14'b11111110110011: Data_out <= 16'hFC39	;
				14'b11111110110100: Data_out <= 16'hFC45	;
				14'b11111110110101: Data_out <= 16'hFC52	;
				14'b11111110110110: Data_out <= 16'hFC5E	;
				14'b11111110110111: Data_out <= 16'hFC6B	;
				14'b11111110111000: Data_out <= 16'hFC77	;
				14'b11111110111001: Data_out <= 16'hFC84	;
				14'b11111110111010: Data_out <= 16'hFC91	;
				14'b11111110111011: Data_out <= 16'hFC9D	;
				14'b11111110111100: Data_out <= 16'hFCAA	;
				14'b11111110111101: Data_out <= 16'hFCB6	;
				14'b11111110111110: Data_out <= 16'hFCC3	;
				14'b11111110111111: Data_out <= 16'hFCCF	;
				14'b11111111000000: Data_out <= 16'hFCDC	;
				14'b11111111000001: Data_out <= 16'hFCE9	;
				14'b11111111000010: Data_out <= 16'hFCF5	;
				14'b11111111000011: Data_out <= 16'hFD02	;
				14'b11111111000100: Data_out <= 16'hFD0E	;
				14'b11111111000101: Data_out <= 16'hFD1B	;
				14'b11111111000110: Data_out <= 16'hFD27	;
				14'b11111111000111: Data_out <= 16'hFD34	;
				14'b11111111001000: Data_out <= 16'hFD40	;
				14'b11111111001001: Data_out <= 16'hFD4D	;
				14'b11111111001010: Data_out <= 16'hFD5A	;
				14'b11111111001011: Data_out <= 16'hFD66	;
				14'b11111111001100: Data_out <= 16'hFD73	;
				14'b11111111001101: Data_out <= 16'hFD7F	;
				14'b11111111001110: Data_out <= 16'hFD8C	;
				14'b11111111001111: Data_out <= 16'hFD98	;
				14'b11111111010000: Data_out <= 16'hFDA5	;
				14'b11111111010001: Data_out <= 16'hFDB2	;
				14'b11111111010010: Data_out <= 16'hFDBE	;
				14'b11111111010011: Data_out <= 16'hFDCB	;
				14'b11111111010100: Data_out <= 16'hFDD7	;
				14'b11111111010101: Data_out <= 16'hFDE4	;
				14'b11111111010110: Data_out <= 16'hFDF0	;
				14'b11111111010111: Data_out <= 16'hFDFD	;
				14'b11111111011000: Data_out <= 16'hFE09	;
				14'b11111111011001: Data_out <= 16'hFE16	;
				14'b11111111011010: Data_out <= 16'hFE23	;
				14'b11111111011011: Data_out <= 16'hFE2F	;
				14'b11111111011100: Data_out <= 16'hFE3C	;
				14'b11111111011101: Data_out <= 16'hFE48	;
				14'b11111111011110: Data_out <= 16'hFE55	;
				14'b11111111011111: Data_out <= 16'hFE61	;
				14'b11111111100000: Data_out <= 16'hFE6E	;
				14'b11111111100001: Data_out <= 16'hFE7B	;
				14'b11111111100010: Data_out <= 16'hFE87	;
				14'b11111111100011: Data_out <= 16'hFE94	;
				14'b11111111100100: Data_out <= 16'hFEA0	;
				14'b11111111100101: Data_out <= 16'hFEAD	;
				14'b11111111100110: Data_out <= 16'hFEB9	;
				14'b11111111100111: Data_out <= 16'hFEC6	;
				14'b11111111101000: Data_out <= 16'hFED3	;
				14'b11111111101001: Data_out <= 16'hFEDF	;
				14'b11111111101010: Data_out <= 16'hFEEC	;
				14'b11111111101011: Data_out <= 16'hFEF8	;
				14'b11111111101100: Data_out <= 16'hFF05	;
				14'b11111111101101: Data_out <= 16'hFF11	;
				14'b11111111101110: Data_out <= 16'hFF1E	;
				14'b11111111101111: Data_out <= 16'hFF2A	;
				14'b11111111110000: Data_out <= 16'hFF37	;
				14'b11111111110001: Data_out <= 16'hFF44	;
				14'b11111111110010: Data_out <= 16'hFF50	;
				14'b11111111110011: Data_out <= 16'hFF5D	;
				14'b11111111110100: Data_out <= 16'hFF69	;
				14'b11111111110101: Data_out <= 16'hFF76	;
				14'b11111111110110: Data_out <= 16'hFF82	;
				14'b11111111110111: Data_out <= 16'hFF8F	;
				14'b11111111111000: Data_out <= 16'hFF9C	;
				14'b11111111111001: Data_out <= 16'hFFA8	;
				14'b11111111111010: Data_out <= 16'hFFB5	;
				14'b11111111111011: Data_out <= 16'hFFC1	;
				14'b11111111111100: Data_out <= 16'hFFCE	;
				14'b11111111111101: Data_out <= 16'hFFDA	;
				14'b11111111111110: Data_out <= 16'hFFE7	;
				14'b11111111111111: Data_out <= 16'hFFF4	;
			endcase
		end
endmodule
						


