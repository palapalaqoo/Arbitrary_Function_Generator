`timescale	1ns/1ps

module	FM_NOT1B(Dout, Din)	;

output	Dout	;
wire	Dout	;

input	Din	;
wire	Din	;


assign	Dout = ~Din	;


endmodule

